XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����c�r��Ż˙�؀��^��J��q��X���*�`�[���ł����1U>B̘�֕¶��>��/�4ǸǡO�&d�Vw��$��Q�U������{�����1�H���2Z#Q���r���i�k�f(FҤ�H�)�v	,�c�����!����,��s/nf�nO�^�����[kҢW�����ۮ�٫5�@�ʓ�1�s�ˎu�+?� R*q�.Sl��id�%:��(��T|Kq2�����m.������z�y+R���k��C��y	��f��y�#��dٻ�^ݲU�r�J\��f��NE\��"a��4�:�аѡ� �֍a7��]��ÐڋN����_����a���酕�TU(�oY=Mv�de椐��o�)L%�^��r�.Bj@��eu�=��.tq�P`g�����mE{�ӧ��Uu_��G�J��m|5�7�(��مZ�K��3MxõOl�FD��?o&7��p�# &��vP6h��s?*���I�g�߼^_g��.���2]�Q�u�Y��x���Q��)�#H0)�Yj��π(���Ě�JR�g�=s,$ct�m���=Hs�y���ٟ�z~�f�wF*���� �z��Sc^~j�y>&n��u=۲�b��ک��+H�Oj]ݗ�+��FFR�Q <����	W�+0nZ�O�ԘuC*Y����lF��������g�c�I���+��&S��;��zVJj��#ڱ��@m��#VoLӒ�֨�����XlxVHYEB    7265    1660�M��a{�n�0i��v�Zi������:x��F@u�gY��2L���?:�]1�/`!j�&���@�>s�TQs��^�0�Ƨ=2�A��o�����
�*�%8�q]TTu�g�Q����|���Y���S�xb�1��2�x���O2x�(�."}����A==����+Cш��-?��מ|��.g*hc�Z�6~vl飤�1״Q�=Qci
"�n�/lH�����Ǆ���z4y�zw�/�p�`�{�l��=���|�Ԯ1"�r��Mf5��n��DҐ/��h�v�t!���ߪ�U'�_�ܴ����UKG�9z�����|�������]�i烈���?�I¡���&����/c!���K�h�/��~�1��\ȡ#)!0��I��64Ґפ�I��TRB��e���|�]F
������V�֒|�,�p	���%��{�ې�=�=�̖�幼>���Ǵہ�Q�	 �^�/X�#c�LQ�S(�!9��C9���b�G�m9��'{n�z���q��]�<���5�YB����Q �W:��e����K;������%��N�GG�c������F�&>%�m$O�S�ek���PY�;Q��}M���0�<��#�r������W?;���6r������Ш=�a��E���Q���2D�� �u�BRG��~>���G�7)țPe>���e�ۏf��g���m6��r�Ds��[l�����Bi��Du���b�|#*�`@N�0Lhv�5�v��k\��y�rDi������Wq�>x-[�a�W�di� ���jd���4���$+�&�MT�1!��I�P6�izx,�$����a���`�#W�.I3uZ_u����t���F\�~~��%��9�)�;7�(�䝀k��g
� T&g/�	��p&�3����P��L][�د�=���}��]�i58^�:Et �>���y����(�
�by����NZ#P��jU�6F��d�BD����خ���:��,�'�G�����g	1��	<�CΧ��R��`K���>��0�]�V�"�j��*��gf�U�*A���n(m.��x��U��R˚��	k/�My�N烄�$�~J�2�66ױ%��+w��ZNzl^�_�t���K��C/�FT%��}/"�%�����cĜ���}s/�z�s�9c�;3�I�c��ل.=�6�isGA��0�a!w���C�R�*��ʲ,��t�,���]!f�*G��w�%�u������M�}5{q��fU	�c1�01�@Ý�U�K�'���/�b�ڷi����>�{�y����6Q%}�t����ֆ� �/�æ��p?6�l�V��hu��L�8�x�OW����	�S��U2���e91%��zAYۓ�� f$���Cq���V�����S΢yGI���n�#w����u�?�W�Dx�u��,1��k���~�6hu�~�H:�t� �bд������]9�DH]����)�K�R�?jH4\�$�Z��ז+��)�����_\���c�#Ӿ:����d��}�)~o�wҒ�VA<��7�y��r֥g���w�����Ū�0:z��p��3�З�p�A;�}���h/�?W�m�	�;7��Ī8v>�� �����L��;�>jJ�M�U
��˄�a�H/����K�}Էǘr�1%��K����_ y���MF�8�����r�/+H�Z�K���i�d��ƔO�!�����6���.��cR������:�5�����=CLB���Q}�B&����>�2�/�pjh0r/ry���*�;��S����:�/��3m�??H��E��wX��P��a�}�ޓ��;߄�+�@	v��Y���<����b]˭)�.�+����v?��M19�<���k�vC��%�d��a�Q8���!�ٳ;�3A����b��S��ݥ��D�1P��	Ġ��.s��ֱ����@K��'���İ��ڠy��񯄽SG0+����1��ɩ��Rg�o��*�NϭZ>äԹ�*E��Di� ��G�����7�:<���=9�-��k��@���N��=�@�&B5f�i�A!�r,�9�3�*p�_<=d���E:ME�4�� ݐ�2�\�/+�\	=���+|��g���j(��/�8jpYu��h���)�F��h�\O��_��p��r���o����l\�K���*>q>��vZlr��\����r
m}����?n�v�Q�����-�8HJ�p�̥���a!u��~�Y&��D͐���Aw_��f�Ԁ۠?x��"(�a@t}�̥2}Z��4�7�Q��N�0,�d͕̈́����I�)�'�a��.�+�F~!4X%�o έw\2s;ѯ�u�<#6�rw��Ra=�G3����7����p���N��7ΖM��}%��!G��ـz�b�?.��7y`��� �	l��%��+Ҫ��l��t�ʏZM�����Oꦅ#�^UTa�j��q���d���{aې�ܦL�5ȗ��h��Ҟǆ!Y¿Jd�\�����sڊ�1U��eZK� ��v��#��pk�ںٌ���H��̭�7i�{�Z���,B1��w�(�jk��8���G�c�8R�I�dSU��B�8\8�ܐ��w�wI����,|�'A�ڵ�9���-��d�����k'��󦭸ڼ0�3��w9��M������D6�r=Z{��9��E���.3����lZp��74��P&���j�A(�xЍ#ɵ��@�3ד1��X�DP�&�Ejf��������Щ��{�rv���_�)�2���#���57�[�싿3b������z����g;���f	eI�z��-x�*�!�gr���1��u�����F~6�w|��u3w�HBb�L/�3�&�j��G�c�� ��n@\CNz���hox�=��VF�A��`i^���V�]�;��{�m$����:����K���c��唜�5���j	�O�M>�$����K��w@@���Y4�����8��8�Pz���}Ӹk&U;�h�����a[(F��?����e�؍F�p�U���<��dY�zj)���Q����+q����L����������;�4����(����l�ӊ�b+���2�ֶ{c.�	e
��uHB}7{_{Spy3e�Dö4��<6�o�w��~�Y�_/Dr�HF�A�K��͜y�J��cl�؇v-~���.�J������G]��S�!����iD�"��Ʉ�{���h��zWI�a�Jeډ�fJ�٥�����&t��ɣq�Yf�Ѡi��!�1���b�)Fh�,BK�U��dl��I'�A��F�[�6��]M�>4@��X�/����_�ɧ�EP�$�'��']X�RL`Fz:��{P���U�7�Mg�o������Sϊ�7�S��8��e�Co�3��7�A�V/:��C5L��d��N1E���F��[�� ��<��0q���1��lk�x^	����rM<O�t��U���,��N.���h%��@�Y���'���K��� �B�a5��NQ����l�Dէ8��Y�_c�v�Pl��Oܮm׻+�� 5 :4��R[F��\�.	/�V;G�+՝��qB�L��$�ohe4��3)T�/O�~�Ҵ:�F�ȯOJ�/��fL���~؟|���l^�;�,��)J��x}�f��y��M�o���>��:�S@8�U_?m���j���X�B����=1|f�ǧ�Ѷ<"��*�xq���3-nꑿ�.�U����H�@nϻx8�QLg,�;�0Z���G<�É��YJ�3\���_Aj�6{���Ԕ``I��y!��0vM�ReUTmN]��ڸm��lS�CS�P#�Q�(�0s���x��A2�6xOy�~L#¯`G�<Z��ɬkb�mR��)c��x�$�#0"@�[^y�J��%�v�-f7ِ���S�3��\��&R�2�`Y�g`������K�e�o�LMZ[���Hʯ���2��V��Ih,����Y�� �51[�<�B1[�9-�?�6���/���^��҅�����Iy��1�G>�g�
�@D��3׽�oyg��K��%@.A^t9�p:`���%2>[$r;���Ip���N�E��S'�T����Kx�!޷���6jg��(zL�n,�l��x��lQ����W�4����u�2`R���g�ꃬ�Ut�p)�H;�=i>�a:b ��*�� �MQ�خČ9����<R�(������:'��'P[��I����/j(�����j@���� (����(m��,��_�C<�h��� m��o��1t�s��;��Z�KP��D�I��۔���=�i��:;�]|���w���(o��=�������@�LC�m$���RuP,L��*0���wGy�t�6�tg�Ǖ�.�o/-���/�m ad	|�4�2�8o��;�qnb��B�{U�X�9͘z�B�2{�;�S�QV�_S}�F�[�/�'�BSBUZs��j���:�T��
ۤt(��Mc[ ������h��z���`UP>o�nl�r.�ɭ(Q�IPH�O;�hu���pM�ܕ�N�LT-�-�m�?��b�S�Q�-Q�z��h����g2�Q�|�j�L(_���`��,���z��+���I���/�vWD�<�~i�(����x y�/���M?��ic@N�=q$��Q���L|��L��$�D�|Tj=NraS�T��3m�G�*S��!�]��s��{�xF�*�zp�T4*�i�ai}
�D^�|���U+"��U&8�6�̏pr�jD�hZ�3�
#�:�6&Ef��(gv��c��Ⱦ��>��%/�[��'~_���%��3���@��k�χ��L�O�/�+h;�ށ�|��\xI[E�4�wfY�����+�����Ⱥ��)�ݢ������~����2�qUw$kO���a�g�l�p��c�k��Ȏd�W��(�k�J,���JdzpGC\Ɓp��2�����_��O$�<#�z��Р��A�#鲿j��k��-�gP:��`�?��9�%>b^��C�8[���B�r���Wj���z�w�=������Az>�yPF����NZ,۠+u��c,�5&�� �f��+��"��SӢ1��2�p9��F��Q�z?�J�����s��h$���ȗQ�ɖ��oZ'�6k4'kB���t@jw��#�6]���x��h��r�	1,��ᓽ��/��z����LV5�lx�I`�Tb�P1݉0��1k��I~N�=c�a�XI�@vko"���<U�������H�?@��&G��K��i���
�Yc�	���*����΄������f}4sʊS�Lt(���;jS+�ߜ��])�A���r�p�j aX����J���+/�:��s�F>�bs|�{��r_�R�4�n��(���9��z|oV!�g�Vbu��I�{@��>I��7Q�,��@���j�rDe�� ��U�-�|("��gm�X=:G,a���U��° Ɖ�R9J���qE@�l��¿V����R�S 'H҉�_,��{W�j�	�X-��0�%9
6	�����+3���gڣ�f|@��ʹx��!y�K� 4��2���@N6@���7�9�ho�E%Yp9�vS