XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��j�����@��C�9?�,d�YTN(F�eIP~%��9 S���{٨���4�0
���₈��b���K��#���������\���I@�A8��o��1��I��,����3RKp��С�Ǜ��h�؟�����3%�.J�d�<%�l��d!��e�n]��R��)i}�5m�<:�w��
����:�w7���JA��ʚ�ɻo���[|R�\���9�%\��#B�&V��v�D��-�Anyza 4�rɶ��O@�F�G�꼛k�4�~)$��1ɸ�d�Kw\[*?6��=ɵ�15!z8$"�L�te.�6�/R�-�X76�M�C����/��"j��>Y"y�ga�l��Z�"�?s��[�����z
J矎B�9�2I�W����b�n����8���-���F�ߠ��W1��v������z��`)�P����*��`���Z�.R9�{����ۛ���O@�  �4 X.�!y	��g��Z�~��3-�p��j�B��9Nڍ ����pQ�Y�ߧ*�|�#�;�j�/N��j+$ȣᾞGk�ה�v�yf!3,�k�B��8��lz8��)7�����2�8qX����UJ?=�����UNf����%H�
y}ewy��M�Ϋ�4 hq<f?]�	տ;a��.	2��U���s@*��KL�#��������N`���Bc��4N��z�O���C�e5�b���>xj�b��?�!��|V��m+{���-�XlxVHYEB    5866    1100���X��#�hE��Ȁ�L���pb��a�#�/�����"�(��F��rC3*;.�r,L�*&ĺ���C
�X��I.�o�e�Zb���Fo����D�#EĘlVY����;+�_*N�xT����5�qB���_9����q��3��. ��*�2�h����
�f���Z}���d�x�O�[�X�Lк��zg[�;2U��.M-�ir�n�bb����R ����b����~��$s�Vc��9/32 �xq�C�u O��[��4���x١ܰ1M;�����W�`0�ыCuϭ  :�#~Ӌo��H��N_��e��LA9^Ctnՠ*�.̍vv-�Smui1 �W�X�+k%�*���)$�|+.�� x�m=ϥ�$�D��<�يs_�ʙ)��yH[��
�$����4Ƣ��u�s���클�%��Qҽ��Jѻf��Z�o��Q�Q�?PF]��M(>�����������SԒ�������FsQ֨?g�on��tf-�h�SY)�.kh�ʹo&B��x=d��&�H��(��XyG�t�*�]�NHSV3��l5��ש��y���'�(bv#���$-�7�����Y�t���=�Î~]�3Wc�ƹN�j4-N�d:�������ʧ��X���A�҇����	��`*q���{������=,��x�&qHgY��+I.4�*NV��
��U���?��۫���-���ڲn��߸�<;Of[*����5EN�iİ���5P�4e$F8/������OtF0�g��vz�]5  �Wy]g�dQ>Z_>�JW:�c�PJ�#~�)%T�{��њ+�_���)^Eg��u��\XR*���@ϩfɞ� ��G�mʶ�)[��6�a����;��&ٺ���GV) q�w:��&iFaD,�u.�EE�����>���t��61'{jA���U<]�)�pF��RT�o�~Jn߳0�dA��k]c�Ʒ^Wf�����3L�$C���_2��g��K�$6y׃����C_��6el� M_��d��5C;R�^ʝ���P	�r'�<����s9��sHlw���)W3��E7��fQƊ�c�����|{�50aH�!Z_}[�V�u��e��o�FE������q�՛�;��L��������}�aO����m�ؑ#�Q2	���|e�|`��e�'�̠v�#�JwU�ig;���B�p?~1��>���Q�ˆ���T����W
Z�M���%ڱ�*�~k���{�41�m؊TJj�Wd���d�̎��N]@�
�̦%��p���;�H���s\pݹoT��LU�Q�����O��q[�~BG'�����)POi,���лx���!C$`��..��O S���q���n��9P�rߢ�'Г���0Oֱ7�8�.C8�� �!?V����;��M��1vN�y�YE�|�SD�.u'�4}�k���|���[ԕ��1����`�O��VV�G%�X��y�2O�۰����H`���qj����p����n�:�Vxn#K�-/63�5Fs�R<��?�Xڬ+p��tUF�F�X��w����L�?�JB�r�=H�hnq��l��lD�{�^}�MpN��6{��bo�C	?b@�s�Y�xC�+?$�d����d}����1jy��r��aR�!��HۛA��B��9ǡ+������{�	`��2��H�'�$���]����"G㻪�&�X?��K�G��+���X7
*�4<��2�_�|��3N�r0KӉ�$%l����4���.Tl�	0$Z��=�#4=�M�¨�C�?qߺ�@��:���,'}Z�� ��#��þ|�!�g�C�VWP��G0v��@w��g�a�Q�������-��sX��S�[��	�ͥ���q�\�#�C,z�oD*�DAd,7kW�	��m~�̛��r�A���`0z5�t�*1�*8�{V��o"�B+��Y?�{u�܅�i�T����c��֢q����2�AZ�I}�I�Y�ޢa6�Ed�jYI����G�"���\ E�@�� <���E3W�V+�rb�z���O�8���v&gR�z@�S�^r�ۅ���a��kR�_2h#��V��T{�"��*e�8#]]؏O� ��j��_������M{H�����)����{��R�������������v�;F�����"�¾�)v#���>I���8%��V�v����\����w`���,�K@eh��"�r(�{~w�Ҕ���C?�[���uK�uˡ�$��-��K7��� ��5L_���\�4�&A���t�!]/.�������\b�zb8dsB^]��+֞Դ�`PW�2���Bu�i����ٗ�2��öb�.+R!��������]���{�xE�C���e�I
��'��]����{	m�P3s�rԾ%��F%���ĕ����V���-���P������R��E��]p��2�0�	"�]�OtI���'��i���^7^Nn���?��߈_LA#���ꈲ�*""��1�<�%�v�a�̛s�Ր�'w؎7Z��ǧ[#OY���`����*��ݨ1�d}��-��!�K��ϰ�'Û`)G8{��e�=t��eb�(V�?�c��^���D/���T%��Cz/�����_O���i�@�k���=����*�ʭR<*�7d���v���ۻYo��l��r=�u�2��kH�6�FФ��M�ӫ��"N�H��:٩��ކK��Iخ/�e	�A;��ݛJ�[�b��ߩ�gی�����x�ަ.z�����XTU�!.�� ��!��[�l�K���[%3	��cl,cs_ Ol�m����4�v�T����O�'�K�1��)���%�F��ѵP�JO������Ő`�Ťز�"ҡ>Iۡ��!=��2��&z[�'���*�r�B�P8|��X��!�w8n1��!��p/���K*�m���z�������������5A>W��3�%n�t�ܥxu�%�H������k���7Y1 d�R^���>�|ž3u��7��ﰽ��5/q�r� J��Øz!��}�@�N|�q�� �zs����*s��Ab��:+- P��.�8�ud�����v�Z�.`d,:ܨ�d��
&	�u>�zd���Tv>��Z�]�߃�F�E7�l��S�����I�U�u�����a���:O�*�]�'���ݟ�6*�}N`��~�7Ԭ����^���1����������2>�#{:�>�G�E�/�{F{d���|�겴NV�Ǿpm�{Z��ߩrι똅����ON�2S$W�M_C�*��W�B�c�+����(~p�;O���ıՆ���W]G��7�;i�$�m�1w�
3 ���y,�?���T�����`�+W�Lw�x��7`hA�8P���I*,��}^�ń��4�9D�F���j.�om�Kԕo�~�>O#�N|k�X�4�!��9y$��A0�6��ҽP=q�ljjK(�1BŲ��Ol��G�.�6J6,,��'O��+�O0:�/��weB0o�SkW����$y6+{C��8+iz��I�l�'?]�D��(V�?hn�ĆKM��+�0&��_axR�,a�!��j���j��N95�
g�;GwVD�'2�O�Ҥ����P�Ԩ�� <�'zSG��L?�RAb��1�?uA)g��T3R+~�j8��|�"{���J�ah/�R���#�M������
�K/W��<+��wN�� ^>3RO ��L�t�N�y/�hΕ�4	9/�@�k,��X�f�w�S)����q.��+��|zH�_d��$����(.e��Nr����4�{$����VS��pb ��k����an#]��i]�*�����|�PIx'a�|�M�y��;�;:`dp.Qͺ��g�,���]�ӽ"&���L��m�G"�Rn@V��v3�]o��Bá�_�mcb%����cJ�����ۺ���Չ�Hg˫U3��@��);��^m22�ŚG��{*�_��h��7>O
�J�|����B���ǒ|��}�dY���*����͛�N|�ʌ\�Z��6�h��8����툒X�L�>�Z��_>���'��l��es�e���Q�$Flp�ש�#�1�ra�����Ja�A�Cn[�J��6שK}�����ά��s��j��O��gE��Bzj�ñ�h ߑ6��+�����л���]��~�p�N?ƫ��a�%�B���{�o��z|7�eS�*M�)����'3�|����{�g��gz�[��en/<h��{.\R�^�Tw