XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Kec�����0�.��D{ʬK��jc��]�Lד�f���h���VBy$ ]���\L|RcY�"��ڔ�Ln��D�T�P7;�HӸ�!�3
bi�&}.Ө���R���f�~5kv���,�����]P.:�j�ȩW�y��(W5ؽ�S�U)Ѩ�G@���9�h(���'w?��&[x?�%�.�����q��e������(�ۀ��Yr�jP)Ҫm�V��z�gl��0�I�M}�R�����ŉ�l�v�}�m�Q��p��2FKQQc4�һ&�k�[��铴J�u��UA�j]�²�9]}�(�/�ɸt;����	�xKޜ�V�v�/-�g�-b��
�8~��囘�F ��P>��\m�R����!O 2Ɣ�KQ���}�b���^VD�uC�D�*C�������/�"�m�	�����y �:G���tɻ�F�g�10��3�L {��CEe�a�y������uE{K�F(��W�:�����]"E�Ӄ3�^T��ɀr2�4�M��>����w�18�nso�;����ڻ^�=�[.�`Xp �̪
I0��Ԅ��F���E+�
� ��e#"!H�˟ǿ�Af�"F�� �$\�%�i�zV�3z�~$�ڛQ5YC��(�Q{^�d�2U�/���z�y9X���,��C�n�3�7��UQȈÍ�Mj��)Rk�1�ĩD=��0���rɼa�1�?0չt�wB-���U�)�y	�Z��hɯUq�si���0��qԊ�p�W\u�XlxVHYEB    1a2e     8b0\��OͲnWt�Y-���V�z�<_�|�Fp=6��	���F�K���_�錸#�]h蚧V������%��\{�Ƌ'X�̩�9;��}�����v/�r=�&+.�M���}�ډ�v�yn�9����{ap��[�,{f~�Y��xpR;_���Q��p���
����U0�mG=)�S��$�M@�����mg$}�S��uE]��۪2��!?N��8�5�R����5E�������c�5.�c[����*@�"�i;dF́x�Ό1A��1����I�Z��nt�
�R���	�N�R0�"������W�5�����#���B�SS���w|6JT�6��#�����?,{:q(���H�y+�̠�B���p8b��-*�\��u\*������L�`taZd�����@Iރ:����qu�p������Aʜ��!K�+��
KF�e�	�(�M�cyt� Z����i��*�ԈU�]��GYF�]��Z��0�e�M�˰�-u'{���J��VFr}�H�\\�{}\aZ��t��"K�̀t� ��
�;��\�-0��6@kt��%:��#u������������X��ɭ0`Á7��h�O�j�<�t]�b���s��\7�12�]f���>�:?�v� �i�!�L�&te��Ɉ�}U��aTmr�2X�!�lZ�E(�\�U�to~��m��bY��K�n�1��$�g�$vݛh$2<7_@2gݔem]	t��W�t,[<ilqm���BعPZ ��K�רe�#BX.?��nT��2�o�Y����~�#��
�$q{.�d�a�%��v���l�'8c�[j!��cF�v���i��aQ��eq��_s+7��ADb��g�L�E�vOT����3 0F:�	@��� y�a?�~� ��r]!Jl-���vF̫;P���Q�M&�,�zګ�.Y��g|i��.m��u������=	��q�<���Frñ{h��=��=�1�sP�s�'��z}�F��Ì)�[���ղ���Q�*�v"d�^oo(�y�G���EHvW�*���!k%/�/\4�z�GQ��a��lcۍs�'ԫ�X�#�M6/����p�^��)��kx�P
�I��誂Aix�}��@�J����+[�S��~�'Gsg�#�%�?s��LX�� �\�E"�_�qw�� �ڥu���e���;0P�݂LM���@�x�2�NO�v''�u�Jĳ��҂���M��:�V��2x�v[tƯn������H�}s���#6���CW����/�&�w��t�N�O�� �!�6�R7l�ݾ�Jo�����&D�&b(Nd�Fʯo�Ӎ��uF��2V��}���si� U��q��-�xu����A1~��\y�D���� ͕�nN^A��8MX�h{	o����~�g��f��͘�m��K���	P;���tN���i��UΓUw���pη橜�@��;*����˖����J�E�WfV����. S��D�/F"��r� %�_H��|���\����^OG�F�_J�4s�Y����ӂ��-Ѝ6:�Y�O�R�W7Q��}�CCh�Mw�.kh�}�'H�ON�o�_'��V�D���m3�ml�J���� m� a��`�J����MT��\�������>7R��"�X����et�V�c�8wu�i�ύ���!�$%���.�Qԙ�!��|��dw�Sc�\Y��\JR���R*(Uu�ּ;���J�$3�׺�6�����\��gjy�L�DR�4�y��6"���L�9�p`���N��\��_�8�����+\�IcI���W��$)�'E�)%1H��1��[�}MyVͫKg�t<����Ѹ����r,��_
́"�!ˣ�];�sܰP
>y�m��rK���0���8F�p�wR)�lG�A��i
�f����u����:P��5��g�j���yGmi� �a�n�i�|�_��e#��Q٭=��Ka^���mCF�G�$�؟~���ރ�B�ν<P�H"i��f�&�	�����d{.:�@3��$Y����7�699�6��J�=`�Z7:Ui6lp!��	�r�s�%?b��W�c@2���N]�=_[��O�!w�����Lk@O�b#+�l�Wo�g�'�Fqc4�*��H�
)S��Y�1�,T*�I���8�ΦU������c����