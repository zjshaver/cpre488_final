XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��h11�0�8��VTZ6�7�%#���l^�(���H�������Kl��_�@��&��5dj�Kv���Y פ<���/6M�tz�$eJV9{&���ʳs�)��_I+�.��FR<)G?�c��!,�o~ha��1�3-E���'�$g�1|R��`�X�l��GF4[��X��rٻ@�jO�����55� �/���g+�^���u��.#��V��nMԛ���5V*& �a#�-:k2@���+��Wf�9�v:��t7�P�g8�ʿ�m��Q�M�F}8!�$���-x�l����\�o�$|v�ɓ�0�{@��`R?}MT�qԳ��5�[�m�П]�Q�K����4�%@=�1!��An��ʇ���㭊רB(��D� �A�Y����v��!g`a��y�lq1n��ݫ$i8����5�+S��t�uo�Mғ�!�Z`Y>�@�|.�+���h�QK�w6�R@hq�!�\.��w�tVa�:�E�`K�FHz�6���bm 5���Q%{���&�r�L(�ȟ�o��	�Ѵz�,1�w�&����.����9j�5rwE�E��p��� ���U��6�M@ �ב�bk#F>uR]�G6N>S�������]���~(;�0�y�3�"�.�g���ږ5��PC���h� ��ɺi��H^zb��u���8�_K�����g�zzn�1�No�J�K�Y,Q�!��ڬ4��]��1���3���2ͽ�uԇ�[�݃�Ue|<��_h@��ڀfXlxVHYEB    aee7    1ab0�"PV6���U]�c�T��p��٧�V���T�}��]��;�pDh��
?��׊7k�]tZ/��u,~Y�=�u}���@@����`���
�#���åäK��JQ�d�����[��Ip�΂��c�t�j��yՐ�V��a�nx�Ic����a�υ���@nO��>��i�����}��zMj�7�ڗ���4I��R|h� s��On 𮐅����`��A ��ւ���׬`�ho�����HW=�3��"0/�j�|�#���MW~ʑ�b��HtJ.����H�]�ג�~���3��kw�A3��n�Z?�(ž���5�A�'X2�~�Gl)^^�#���mE� J?�i(�^���/@P@P�DW0�x$�E�e��B�dv��H{�cD��L���Rl��^v�jJ0�x����6���)[&Uݬ��>��$WR����5$�P~"�ǝ>[�9�]�L@��X[h���)��XHdnE�B�O���3�2�~K
p���]}�%<w2ż���ʣe��@.�7%���<�!A ���_���:��=.������2�E���)��j�3��\+:�kq�A�\�,�#>�A�u<�������}*�2���t@8j������ߦ���~�����UZ��-���o {����U[7���3�[��U�
zR��`7nW~�h����M� �&�"�r�6!��e{$�/F�C2Y���:�_t�3Ok��oQ@�Kr���d���[�J4v=�=��А��V�/36��x_����;��T����ht���b5@��}��OCG��n������">yغ��wN�&�9�|�XU����#�����΀-\Cw����S���e�^�5���u����[A��70�]�Vqf.������7�>� J_E�Y�=�[�,N
)�Nص���K��[�ir����bnx
�}N5�1�ϳ	L
����6�Mԍ�:�F��\�����z^~���b���8}Y����gs[�h/D����DUN�%r��pHS@p�:_כU��
�')֎4[���/�df�l�t�2H.ڛ�<�c?�91�o��=�))]�u��Oi�=��-�s����\sjy�X�ˀ�%<quÎ".,9�֦��PZ3�㨾s���!	2#�Q��H;�N�!��PI$�{ǧ91�d���`�<)���<:y��x�ց:d�
���msY`?�ےX��@QH䩆	^˺Z��\R��-p9E��%�(���>-�p:h����3;�t���VΙ�\n>��X{�ϝvq�gi ��[0�&HI29C��b2�r��_(}���Fh����yj@�!'�%�u�Bg#�=��%;br*W�2�;�u %�Ȯ��ò��Hό���������AW䙀��j���yc�,�0��ϵvI��/�m[�fI�b��*hL�䔐�%0��^;����.F��5f!��A��ʅX�]`����u֗\*�'��>!�>=��麓������~6�"u"	��CL�&ޔ��=�([���
2Mbx-����	�1�kz#�c~�ZN*���ޣ��S�;�GH���(I���:�_f�:�M�}CӐ�i�B�JJ^�G>�1v��K�À��.C��6Q��>�5�SHj�ڮ��@=�$d'�K�Q4�7UIY����H��F��6zƽv�߷7U���Cy���
CX뢩)۟�$M(u�eMT��T#���K[����f�Jm&�v��_�}ʞ��gM|���]I�gi�0[��k���#�X�9�(ZI�՚MmH���$�cE{=-ߝ��x2�w��찢��N�4�Mc����Ӈ��x�:�iS�!�\��f����zlrN�d܇���`��F��/�h�(�`ɖ[<�)䩚����Rp��	�N�N`�J�ʦ�����Dy�@5�3�y�]�k�8��Ƙ|��3<g%Ui�@�M���Ŵ��uB��\�Pa����7)�~��ޮ���P�v�f�'�ޛ����}�NœJ�3,e�t�V[xL�����N~3-^?�9t͛���7����v��6f����f�H,8���*��S�J�U��z���{洚V����id��ck�xXNe�1����n�!�-��a��8��^�����6i�T��n�j�!V	+��ז�(��Zp���;l o�oIQ�|�������D�����F��]V�Q'�q�P�e������Ӿt"���]���HZ�΃72�����!���>Dn��0���舔=��� ����q),z4�alzS�z1c~u?l�`>_k��H�-��醙�z*,���!4FPu��v>)�iα�-$��� LOj���~��F��b�}��Ġ�q�-�M��:?��q����<݁�f�~/���J�S?���IlG�Gf�ݹ��^�|�v�}MOf]�/�.�\��:�eE���h팂���E�H[e���{�FQ��N�S�p��}����5��P>kpm�MU�(^�׈"�D�<����k-d���Kd&�N�3�+Ո�53{�_�}q\	�~M�&��L���1��	EB܏��W|q�ꙗ&���:�1-�7q�ۖO3���fN����UV+k�Q��3X��E�?���V<��<���fW�&����1�uE,l���c!�bOYY����-SZYE8�;*�C76��g &��@��a� �V�����__�>.��L�Y����q�{6'��bgu�h����$�
	ܨ���wȆ��P1^UT8_$\y��2�\ɺ��
O@�9��Q��s
���cG��y*Ʃ���G`\4u���J�R�E���N�k�k3c��g
6r��`N�樾�dh@�^���%;֓��;���\\�/~��w`���й��e_娔j,"�����Y�~��x>e?XGr�h��m$!���J���V�`۹�U���)	��[�}l�� :�đ�!tXW��S�9�৾l�N��Y��l>�Đ��C[��G4#)����hV��]��[$�/��P8�c�N�K�ԇb3��Ts-���/'�U^����&<�����߰�v��P��$8������ٶc���4Qj1��U����2󓫇�2�	��o�EsV�Ch	3�c��*v�-N$g]X�U����#�`�c���yN�4���*}�������ϹkzBڼ�����Z��e�2��W/���0�?�L8�Dv�����^�	)��u����;i��mh9F��:9�9	�uK�~�\�,�?w�.^�G�ݏ����73'��=�Y;���n%�$+^�����a�)>ڢ�����}d��#�����?������u�3�fI9.�����3�5���,j�"iF6�u$��0���P\`����Ϗ�USBC¦Z���4;�q�:n @ꤙ����x��m��t`#��s��mC��c;�׿DM�k)�F:���z�T����V� >�ى_�����Ƣ��l����>�4�Լf�]$���sUm�(�9p�v��ap7T�S�h��?eO�g |��;�P�a���IDK>��z®�
�g ⪳��m��s���1#�.�R��(��!�4�0�s~7�l�P��	}��هow�G�+t�U5�J�8��[��P��_��.	wd'�cY���D�1�F�M#tfj�x6����r��0��M��a��)��b�<�Im���:B�$���	]��M�΁�G#T��h�?&��:c^�ۆ�c���ov	��nvN׋��ݼ�\Z{�:���wJ������&,��|��|�\ZC���%N�=҅=�9�]î��Iy�>�����5�#C�r�Z^��	��r��C����P��(��U~�2�AU!�uY5�EN���l�6�d��!ʆL�ݚ�%�~�g���u�1Z�#5&J��Vgs��K��x��t�aa
c\�]��<�&`C�:CE�m�|�ks�hg���:9��F�AL��9�nX�x�OCeS,x�}v���V� �:f~�gː���`ͤ����r�Ё]�T]BC�y�j�50~�Vk�SE�6޻�n0�3��.�f?��R�!N�L�gu�ɭ����������l�L���˃G]@;@_N�v�����-�/��"��l���rX�|q�V�˂��$Ψ��R?3!��G(�4iM���S�tf#vޛ�o��v����ʠ�x��	D����v�
l��q�WH�{r�����X�n�dj˺��5�FIe�\o�����twl[��`V3mD_��5$fՊ�YV�=8��f��nR W |�e�Ry�(��8w/&��.��Pz)�e�~�'Q�)$��ܱ���JܜP�Hm(�=r����t���#�T����{Bc��?�8%���UO:�ޭ�3�Q����Q�����/I����2/�W�Y�����<w(��X��m��v'��h&���1I_�1ZH��h�Ҳ�e�{GUx1��s�K��h?^
�]e�,��V��8(*fÂ��X�SO�)�̦R&�!�e�[��彎ke��g�[6O�G���bu~z��~O�e�|B�a�����. �!���س��{�Ĕ�g���^0�,�Vሩ����Ip1��|��{$Ln_	N��sEѫqĽ)@Ϻ�kH�!��ݭ
 {)�����[N�25�]�+�a�T�1`6�9�������z"z�<�z@^�]�Q�%B���e�Cu��`�sj93F��;}qJ�L=X�0���;�np�I~�ř�����G�(��n��]��v�� "qv?[f1���h�Ξ3��P��8����7�{��fR���F�xFm�EUu��R��b��%e���YQ�ӎ�P�U��G��c7R��E�u����7b�(kSa��3�Z>�vN4@�OMk�����*�w܀]�$W@���/9-��ߩ����&����͡Q��pq�
�8"x�o���g.LɻE�|&�Xp��.�3I�����ڲK���5����z�x�>�#W\$цT)�:Ap�e�e&��?OJO����b��7�M/�����
ϛ�JI�ME�eSK�JV&AXb��Z��	Oz9јF������W]/�H���"B������]�A�T���+�����9К�trio�U>.Œ>��дZq�%�>OU��蜂ĮD�߿1��~I�4��	�����5R��s�r�	��m�wT�&;~bȉ�ܩ��#��ɺ��*0�iD38S���^1�D�]�
`]�FVS�{���	�����Td��[ g��W��Jʤ�A�Pc���z�DJ�F@Pukr �V��h?Vu�6�
�C(���|�?1-����g����w�	2�ڝ^��eM�q�#U`Q����[�4���sJ40!�y܂6�c�!�ћY\E�Qh��67�ȓ Ά�C(��m�.�#������☆!�̃�,�{�ڰ�Xw�+�ڨD�y݊��5E;3qN&!ֳ|Ҧ>��*̀��۸{�!z`�*��L��dsS=��<m��&� ����. U�n��fljz�L���O�@��p^֋���Ӫ���W���ʔ7���)�J��5��\J����!W����0hsK�Q�0�n�*a��b�H�Q�Hy��ʉ̖M����.Ǿv2c��xR�il��HNZ4��v�d|iFe(Ud�eY�tȵ3����f.^`O����}�{�30��j�x��W�ޙ՛b���Dp���O�ͲVaP�<��$�mv\s�do%�c�op1�<��%��*Y�Xئ�X�X>
y!�;IŨ�π%f��ah+5+[��D{�	�ŧN�zfU@}��`�����r��Į�&����}�HS�C�� x��(P+b� ��8����#µwC60$�b���YW,�=����`��5�ѳ�H����Z�Y�Q�	�C�0C=4�+7��e��ŘMU
�����d6�:).A��[P)x���Z�j�2��MM6��%�����t�)����i���;�O=҆z������*�v�22.meA�bkV<\�EU�^ ��&���}'_��6oNw��oy^aYĊh���KC�2)1���zR��)�P�Β�%����yQzr�O0���T��Q�v_��U��X��v�$gh�2�_3�,O�3�Ǝ���%�.r�JĶ�?>R��FIT&Bݎ�go{��A*);G{KM?�d���m�����BXŇM8�m[I������sǤ��L�66v���\�z���O�e��,]��jZ�
F�*a+�p� k�+?�>貱k?Ⱦ��~�{�q����	�)��QIr��59�j1����-�+��yK�K
���{�~D֝Ykd�*��W']p��WD��XK�}Y�\"�e�ZN�R��(��S�_�qM���{p/�� �;VI�.���fȺ��0)^��{��.�!iY׌����1����O<V��
�Y�c��s��L s��g��[ ?�af��Y6���IvB�#Ӎ=I��F�':_���t���P��GT3�qR�Ӣ���+~�tWE5#ݑؓ.��OW8�lao��f�7%���˕�;�X��k��Z2''��q�bB��J�9lR񶖅[��	슁	(�ݓg�.��%&����$Y��4N@�8�Y��7x�'�t��D�	h�>�@�[�3C��c����~n��
��BmEZQY���ɮ����j[�;Ss=�êT����?��>�Y߂�?�����ϚO[^��
�0[��Γ,_�|���e".^1�r��N_]hd�"���%�i>