XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���v���!j6@��+��+xL�?��8�t�b+�L�*�L^�Od�j%q̻ŪQ<�ͣ��O������n�~t{���q�q�R�����Y�i@/N��<x@����l'~�A>�$�xG��H}��Y��qXr߮t����t\%H��Nw�9��� /��L!����D����OL�y]"G�K�h�_+wQVv5����B��V[s�ڨ�xT����tؤ�"�$��c
�e8x,���NX�`�J������jAƯ�ow�k��h~:Xx<��j|)��Pd@A����?E[lq�3f);�R oĭض�ׅ\��蓔�!�b�����򲵵����;\������ΐ�����
 �;}����=e�R[O^�B�u�.	<J�������ˏʕ�<�g�d�+�&uM��\���]�zL�C����+�a�$��CI����FS�����SC�468�P_yL��RP�I�M<3�2 h��v���hq��H��^�!�3��7KU3&=�����}��,f�|d�@�f��گ ��<C��#c��xˬ�;��{+)a ��f��9������7��*{��ZA�~}��;�>�\����,[dE����-������"cg0^��jqFNsr/���VΑL��{�Vl�_{�����q�ԭ�TJ6�`�f[s��sw�]9e��>ߊKcsir�Q���@�Tc#����)�$P,��7��'R��������!�		UM=�v%�0���������XlxVHYEB    82c3    1970�E!��8�M4�F���g��?t-u��~ӛ׼);=�n���]:3lDN�����x�Tyx�i���J�G��mJF(��K�����_�H�t�7�	��q�𱬵�[ݡ���[���ߘA�4z<�ps4`��e��
���{N+ ��B�L�a�ά�3_�P�:K�N�7�Y�Te�4��iL��0�J�0�q5�0}�Te��6�4����,��2|w/�=�0�� �|��;>s�+�}���Z���Ís9���Q��϶˧�\4$KG� #wB}��x�{�@�$�|dQ�=���vfS�[?Ɯ�����K�2��g����!s��gU�*s�`~\�7���o���ÃI�Bg��./pޫ��=uqu/^i쐲=� &�]��8�A�h/� ]1K�X2�Ei���+E�3.)�z�R���6��\fd:|5�k1��87*1� 4D�.�遂���ҁD,�9����cyZ�~���;����
=��&dt+��q�G@ɣ	�76�㣳 :�ټ���J���Z��M��28���d�m�~Kϧ�_1_+>|������^X���8B�r��6\�~]��"J���J�a��Q*���EQ�;EOǳ�����r]Yj�8�-�b��g��;�ڀ���T�;��A�w OZlm'��3zmp��m�U	P�u48��.~�B��\�,)�@�g*WvQ���&~m����5Z�4�?,cRY��F�E�ڞ����d�-���.�R����}��pWt^�^��O�H��߰~� R��Y|@S�CRw��PI�����GP�a	��v㧏�[@CL�����2Z�%j���Э���3��GL��D���
��G��
���`A��C�{��2ү�f�h_v�^�^$���ӂY>s�;$����כ��SM���@���RB�.)I��v"K�Ugq/�ϕ.�6�0��k�i^d����s�{��u��6g�� #=�FD;5c�A�/=v������9�b�L��=����d��%�=�$FM��[�྽!f����������T���:�8�؛U�A������}uqؼk��W;�:�W�+"�GK����#��um�*&�L��W�L.��K���H:矢�X""�:hf�'ܝ�l�C�1Y܃Cs`����O�1��^s��C����ct�K�$j��j��Ԓ�
luU�2kT��Y����q���#y��R���������N�_�KIJd��n����4�"�ku+�ncN�8OX�*	)��܌ +�	 �ĲM���l�WAײ$H�t:Q��}qBs�� )6����G\���)]�9���򃖨�`-�m��ݵ���1U��G:ti7ԋ��-��է��w}��+�B�ޓ��B_�*�hE��4$��dzjc��"�12�ǅ>� �"��I�h���+�a`A�F��#�h�aOZy �HEB������1���h����"8Ր�H;����xG�ȴ��<����ؒ��
G��j<@��E"U�:z)�5�Ř߲g]��7O���en� *�(Z�	 �Dd%���6�G��e5�&1��]���`�O�W"�ZO�v�+.����������ߋ�+d����(�q���ذ�L�y�d�Kǋ>�|�"f���]�a5�z"x������)4�\�ǽ� e�Үq��� �����Ƙ*��57x��o�]�2���mZ�_��_):,'I/�>zlz���tR1�~���B֮�}~-�xs"����1)��
�v�Wހ
�"�^8�}�����UM�f��
`O>y��p�Oj�#�|�ޒ<��cDw�u��*��+aw�>t�!D�>�)���"�"�
_[��e)�ւ�2�F`a`8�Z�3	��	�sf�H� �K<0�D"�.���}�g�Գ�h���,l�GZ+�H"30�}V�VY;#��\�L�VN^�c!>�e) ���6]��"�VY�S�r��w�y����30 �ɐ'@ߛ�?�g��,Hk�����3p1��9A�פw���Va�����s��j%���ֵv��B����o�y��"���e�`넋��f����L�b
�	N�8m�+�؁���!��֪L�zک�a�?��Ě7�Z[H�^Pڽ���ĥ��6N���&�����N}h���z��_��	 hZ�)(�	�q;�,c�L�MA��k�b�44�0t�&¢�����+�D=Ұӻm�S�=�����M���Y3��#L��4;�n�$�i���(�߹Ԁ�MR�˷t>�N��>��w���M3!�F�4��f�_�yer��3o%�p�j$x������f�f��l1)D���洖���'\�
�W��Ӣ���
��i6���/y�v����Ժ^VB��Gkl3����)�w�C3/��#���y��_v"��tjY�.�>߸������Vtz�vĤ���_C��#>�`v	��S4�SɄiZO�� ��@Q??T���q�ވ�yv��5�
�Ρ-���@�л�#s�D,�rw��T�*������4�Be�G�~	�↢�UQ�4U���DӤM�׽~G9�>�|�6^܋[��M��4���+�)�M3�uD��93�N�n�r�s2�����ޑ��ԶZ�����S�=Ro���*��h��`V����G����~��цD_��ؕ��~�[�U�$#	�9{�N16� \;)�S=֛Š�0��b(=�x	�����a��o�޿c�nw%�ˇs��i�<��g�����ME�!ܴ���K��*�*^[�+���dM�X��us��~�!p��� �0Y2��Qo��K�����K�����>��2O��O5�Ņ�rM�F��,iI�`�Ov�2�/
7�~�M�R�<ŗn�З1W�����£����s��,��)�l����S������e�υ
Fd�*)`ZڳG'q��2J�����(ݽ�\��_`/N��J�@��9p��O?����S:�y���GO�/9��ݜ⩻�Z��G!�)�0����I�u�����y�B�y�
6�}�S������u�bNs������X�.I}�<xf�� ǫ�n�"ƻQ9�*�W��Gm���]1���N�\�<�
R7��ԗt�/L"F����cS�D;y/�K����z5;s�����܈ð
��Ϧ\�r��a�z�A| <ր���� >��7�'iR	���v� ��+[EM�Pع�7��T�c���iS��<I6�c�D�2z���M���tlX��u�2�(rpVP�<���qѧ��K�"�:ô�BJկ�=����Z�i;�b.S�jݱ�S�,���{fp;�<ݙ����%]+�M硪�x��X�uZ�8#f�qv�M���*��_Ŧ9���<u�>]\�ϑ����;��ݴ7�2�Qhp���J���".FT��3l�K��.�S�� �����K� ��n��ޝd�P}��U��R��Qs�? ]�s9�W�+�/s\�k��EJ��=:%���V�˹3��qK���kޛBY�qA��˴�Q�y�I����]��oΘb���fZ�'��\����!���p�0>ԕ��8����2c��	"6.m�@�x3�伦��:^-�$_��R��v�Ў������3�����J��ˢ���8�'�;%*�-��G��MyrA?���A���N������c,��"(�G�>!�d���	k��
1I��o�*���c�˝����wG/���l�8-q�kQ�~����2-<�G[�MO�(g���}! Z!�g����x��R�PHJ��E�~�ܮ������Y(t�8���[� i��&+
s~�t�$b�륐�G�(��{��^���$�G���u���0Q����S5 D9�kv�=_�1�[���2y�crwMKlY*��_(�
9�B�Ԝ���һ��p%���� R�
.ʮ�5��}\~V�0U���`%�3����_{�8����/���
�  ���qe�����+�����C�8aN�_��X�u.�(]�TE��x��w�NZ�����"4LΛ��mX�DZu�s�s8�.��栤�W���=�m��i�/9�%�̣0�V�.�<X�oIy����Ʋ�Ni����3�Hy0�Yv��i�`��ȏA�b��c�� �YfY�ݔ��t��<:�@��F��������VP`Meb�fY�Xߡ�︗w�3_��Ő'�ԗC�$ԓ��S�h4��@��\��k�j���6��A�=tީ���+� `gQ��C=jh�{v7���d�q��h�?S�a��j)�
�w�^��^d����ws����`m`�l�z9yʙ�җcͪ�%��ΰ\�^��ˍNU`, [B�=���W� g>��s�])��b����9�H'DGE�<�!л��x5k�����%s�r�4gc|H��d���o1:�������%�«�IO�$�V��X��	n��@gP�Ji��s#�lF�q:DI�9�Bm�x���q���Vf{,4]r7�*$b�sg�eUV�2�$��,N�Da�QG8��v����.s��ON��J��T�͟nAi��|����:	��"�5�y@ʓ�*�U���X��4���0���skl�#���Ȳ ق`>�E��}��w���ܛ�R��cN���Cg��	��<����lD�X{�Y����'�5�#�S�^�V���1��5K��uN�,�CQ�\(&��*ا��
7$���t�p�x�M�@3��aá��`.�j����&$�G�/�8W�b���qU�8H1��z;�qҿ&,\-*��h(�yZ���F1��"���Ԉ��D9�#�}���p��ۮ�;�,)v��e᎐�4��̵xb�T�H����Gb�'����03/�[toI|/��Q�[��.���j�[���vs�G?�i�!ɺ�৩����N�L�H�If�]#�f�R{N�6::����w�]�e��h�Mηj�җ�5z%��)�YDv%���._�;NH�0~稈�{���z�����%�wV� 7$��PС�:�Q[&��Ԩ�� g�G���[W5�ѫ����5��"�vGU�0���X|S=u���xN��F���d�z4zD[����RB��eht�*o .5%��.�$�`=�y��xQ���􏎋"�,��5�>�Kf9��S.مZ-�� &�uAEM}`�:W��%N��/��/fC�%*Y��g"�Y�2�o�%3�F�u�r�՞'t�����_Ǆ\2�3.�*"|E�?m�CoC~q�Sb��$�Y�s 7��I�׊un=g���p�J2����*���p��4.��VYe?K�#c7(YjW�g�9,@�8�zJ��MI_�.4���5���'ˮGM�'�N����ɡ&��tb��� tDt���d����}2����
��K�#d�,�1)��������ɉ�?��M���zJ锻u$y�/D�dǧ�8 �c'����.U�M��SgF:&�LX������0�3�E-�C[T�*�R��3YG�19��Ҁ�~h��8!(�_�tk���	�&�:�ݘ�[b��)�dU)b�	�MA1�a3�OI�%t���no�m�u20V�悱�4�wȬ���9=�r�^��Sð��s�Ç�ϯ��>&��C�H�\�V3���{5�']|�g���Q�Ǣ4��"���܋��W�k�`P,�|��H)��3hA�����a:s�_H�� �������)�.N���'�}ۘ�)r<��e�l/�Wy�m���Z�T+e���[7��/�6���b��m�fm8@F0`.�czKƲ��o�%�a�Umѕ�WLW[K��㚐Ć# ݧ}���Y��ǉb.��0S%0�m�B�U�.�o½�7z�ٜ1�Q��\$�3��m�c@F�u�/�
v�G̀�'��y��t��L��쾛p?�䪚3 �Hd�eHb��޿5�a[ 9ʵ@�c��K���TMo���`!9����7_�S�Dp�7�=�0z� �Cc gj*v��Ҫ#�T�T+��:z�օ����;3��φN������K@��{c�Bo��rg���:�O�2���n����Xcǌ����\ĺ�қ�P##l��|�,���&/0;t?�����,p��Z]�H@80�NWo9�
��i���,�����>�,�DF�r�0�;H=�� )l�^n:
��X��)���9A��k��yŹ���6a��a1}���I���祮�~��ﵭ��`�@����I�{�6�g�@h3 ���&�K�S>�
� [�g�6�9�rB��
.k_�5D��}��9{�qd�t3^�� 4_�V��DV!z��u�[HQ$}���T���_gc�h� ���b����ά|��������nD��h�U$*�wA$�7o�*ӭ^,�R�=�cɛ`�b��J�v�G�x�ӌ�����ŷϮ���L�-Z��ר`A�Mf�)P��8�a�fY��������