XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���==LAe�	��!�=�o)���}�IS
/-�?؇]]�Tƽ��v��fha<����B�ca_j�Q_�r��jz�:|�|&|j+Gc�����]`�J_���o4����tݶa�#(����x$�3|��T�M���h���_Fs��9n�4..��r����+*���[��]`��\�}��}��;�����m���r|ZUA�K�[�J�2�b�Q2%�J���Q��j���#F��1o���ZqE�bu�՜u�Q�q��͓�7�y��_)�,�z�z3���F^*�(���H�(��	5`cI�/���_�����{
,q��ycY�p�#�%��"Jxb&�^܍�P��ⳋ�u)��M{K���:�Ý���:�n�n��$�`�΀ZjO7����F�}�E�)�Йף�W�7>��"���fRa
]sDlk�!D�?^�"��[�Ϙ`���c��E��!���j���˴�*/�s�1�.&*���!V�N1v�!:�����3z�ґ�;�,�`A�cS����Zi$��|L�(
J���4���!J��7(c�Ƚp���ᒣ�%�0�8� ��ԝ9�by�f�CQ��oI���ߗ����M�B�C�s"����5|v��Du>��^4��:�Y/%%���6��׸�
�{X�bpbNs�"�y:��=��	cn���e��Q��,dHb�#��@�Kյ(����x�YR���)b�ڸ�%�a��X8笄�?�&|�Iw�1֑��fD��B����XlxVHYEB    13ba     770�)��m��7�"���j�n��Y�!��iݍ����^-�qĒ�z�1�j@�d�ð�e�2��{�Ͻ<7$
���Q�(|���hd�v���	~��t9[j�MOMBL��f+LL_��bl���Ϛ�"JWE�ױ�딷����nA�VI�
P�8��؈\��W�9j~������c��Np�*��@?�/G�R���eo�>��֎x'����Nӿ�gPlɶ��*.�\x����&oE7)"�܀�'�4�L@t���zEƛSn��,
�sv�S�*�Q�����-��4�4/%]�1�Ļ���u�8�����T�`�i�/SS�G�Y����<�G>��k;uJC��z)Y�/�0�\��!�V�A�J�?aD�������;�&HVt�\/*
�A�vQ���?��pR��ɒI�Τ��D����V��]�.ʺ�=��2JS�ZE�n�B�O]�RK1r��M���'�E��U�SdP{!~JdVox檼U9)8n�S��P{����f;a�SVkK���hH�>؈2^�dC���c#�޽�|��6&k�Am�>l%��C�L�HB��F�Xjn�^��x�7K9�H�}����o(J+�}�u%pU�7&a���]J{Q�f���΅9�|�u����7C���'�:�zY�`v}$�?曘�I�@Ɩ��mBz��t��lC8!�n�s�}��*���'�:i�u�y(s_�;<j�jHմ�����?�w3���=8������p�� ���P�s�=	�&��l�S�Q���Q�����+�H ��YR-��Ʌ�_���E�-
��a���K�������$	�g-���������^�f�KM����¥30c"�W2ζ@]������uD��G�x�q��|�e���(D�E��\)U���{��·�����������C ]�p��-08�����z�N�W�������pA�rv[��Ir�Tۛ^��f � h�|�+e��v����ąj������n��Hu�EY�a�3��D����Bȁ �s��l4�B��5�O}
�����Nw�ؤ]�|4��
��
�,��� 뇬BK �łA��II��kcԱJ��͒��	=K���#�f����'�����
uW��X'�Vw��L^8'ϛB�yt��a`)h"�j 
Kԫ�Ж��o�MŇ�u�C׋�m�_�����cAe��pR�r��:��6;��=�QD]+��<�HUg)����d�H���':���`��� �h퟾��>�=�%",�;e8<�bܼ��69[����p���0�<8k�/���}��=n8�D�V�c=���$�m��-�Kl�H�f�����.� �to�ח*�E��h!�p�����P��)l��Q�vY��7:i��1�'O]�I�����㿪ۼ��Gp1acxw���q���������Ə�bf�PNqB镼�~�o��;/�G�&fE9 B܌A����A�|�e}٤��d���[y�2�U�Z�4��I?ʏ^�d�\�<fTnj0!=(7L0��ܖѱT��/��.�%�򻕠�ZUvl�?d��J��?��lX�R��ih�X@=����R�Z��F�^�C6�X��c�b�q'T0e��]�Ӈ��V	b,l����#W��*��B��\
":k�߰���dWf�G����k#W]o!Ŧ� �Z/�DW��jo����ħT��l6�U�3:�����K�܇�>P��Z��&�|2�"1�l���Ud>���v�p�޼�����U����3>C�0ˋݽ������iO�}��^\��Q}������vZ�ݻ��$��(�ĥ��8�		 ��!�J/O1�������er��[:x������>8Vk<�� B�k��m<߮(��