XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��`s���9^��b)p+cT���~nW�[V+�5:��l�`�5;n~��3��S6�2�������y�Hq� Pґ"O�z��!x�V�r���a[�R���k��8e��&���c�8��H�9��[�P˔m�`0PY׿I�
��09�S���PFd*B�J�!�S�~�ﺘE�y��p,�!�z����y���Nf���mЉ��~a1��HJS�:3�I�����'�HJ��+�ӛ�F�A3$bK�Kf�g��i|)�fj�WCR��E�{"I�0��J˧�	(�~N8�b<l����f��*j�+A��?'z�$��};Pj'�4JW8k
� ����]��]s����e�����h&N)��_B6�{P�3��-EM'x�qa�<�7돧x�u�0�`����������ĸ#�3��h�=��&��GFW:h������9���?���~A����آ�O"��|��S`�:��#��ƝR�����]1/�E4�v����*^�~P U��TX��{���1���]�Ü���F,M�N�W=��H��5�[Z/O����ii���.^6	+�<`CFT��Y�:�u�H�M:��B�S���|f���h�ąj:��Wh�w���ng t�-��~2!Ӹu;Wt��qZ�@�ܒ[�Dh{�nb��D����PD@/x��;����h��3_�����Հ��RӺ�:.�I|�On�q3���$��>������z
�-�$H,���3:/��tXlxVHYEB    1421     7a0�(S���ټ���R:���
�.��u�ϴD�}��-��m�_��:�Ly�x����ﵨ>���r�0�e���q�B2��Q��w��Y�(?��NP$^O_�r�����"1 �������i��W�Q;��o;�a�>� �]���{_Ags����)p�iɥpIzc	����DI^�6���9�:�}F �ӊ� y��6PΗ�ܥ͵݅ۺFik�T�����?)�4�û��I���=ݖKX�4h֙#f(���mU��n$8�3�IY#��á�ww� յ���0I� ]�����(Ąن>{�B�\=�}~���P�a�6���4D�I�l�5�(�	#��n?������U�49š3��I�l��J��!��z Wh���� *b���YD�.�%��iЊ���O���ȟ�o�s�r�D�*kO\4��<��eD8B,o~�W���G/�t5o�D�.�c����a�?F���`Η�"?���F/�h|�>8�g�I*��1� n���X�_�,C�1�I��{V]vo�e���-R;[ E�Ch+g��V���Gn��t���]c�;c��r���e��O2*����	��M����t�e�9
��	j�ΕI"o�$�����b���%�,��5}g�D�a��!��z�Wɾ�*1�$��7�.gԔ�U�\ٺ��޸2�2fr#_\oFsU�a��ڛ ��?���'����ze����+�$#�q�Fuo_�sL	=���}����0������_���I�����S����#�)tB*m���
ُ�(� 's-�>+��q�o����ùH����ji��o���ժ.d�����էu�jS�z�<��w'�4W�񅯋�%ԃ #ھ�Q���˛u>~1���x���d���Lq�����Ҏ��&ϖ�M�?���Y���'��T��_�6Lx�ƹ�,�-��-��Ě�R�#
�Xc�p��tZӽ���.��E�tl�F��y���s���kC�\���=��M!�����0@F�I��f���!x��/�����È=�n����L>�a�q�xp���i�b� �$���I�n���]m���=���z�S|��o���ӝ�
WF�)��)��@lO��8�c%�a"i!����C��̭�/�ׄ�E�B�w�#���d��xvL��*��ن�z�����M����E��F�N�;�v����X�砿1]hX��:�Bc�h�O��#S�G�j�֣�`� ]d����M���H�.��3�/UH1@���)���A�?�&X�*�o�Թ��K�k/��C7�UC�8��^��|�RF g�;�:l��1m,�n��=v�6IC�Qn���UoMc��-�E1.��#���u�v�&Z+��0��j�>OЕM"�'��3�0�fl#Q5�
a�?r�!��;�e��n%/���^o\�%���ª ���%@g�q��[���XK�a�$� ���q�|�|/!P�G��xv;<���Y��#[f�97w}��i��y�@[� gE��pg�Zk�;��� /l�A}��K<�X��rz-:5�R�����Z
��8�R��̶��� dP�[��HME������}W��F�j�v:"u0���E_�	_��IH[�FP6�l*@x�S=�!
�I:�vb�c3Xy�G�c�#v����z�[��@��,v�0�yg�`��cZe执_�]�S����t�`�:%.Q�=�>P�C��K	<��q8ۚ�h4����(�w�gTw�E"3�v@�{[e[�WQ�r s2�BF�)����K �`։��m����<�?�.V�d�~��q��'|����Z��������$���o�����#'W!RS�pﭰ�%�AU���m$W�ȿy���4g3-�,�^�c�5�u