XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ֱ$��3`y�T��dV�	L>tb����P�{�H�Y��i�G-(H$_C )"���8�uՌ�h��l�(d�{�vyq9�,*�f�+
�ɤ:6��wZ�-q3�5���Q�d"��ۍ��~�\�B��P(n��xX�a�H��f!��S������7}��Kŧ�&dc^Q�MɁ6�Tx��j �N"�#Nh&i��\�c�
0� {�>��@�k�+q},Uoe�׍͕jb�jh�<�1e�M��D���UqbP�-^�@��:�+uQ	P�S��嗁���䏓aH1J��!�]`�LJ��S���""} ��A?@�� W�,�p�I����p� ����;�9�I^���p^�����W��f����t��I~�ϰ���[�Ð�C����HpE�-��B>L�:��]o����'�����9��z�w�R�m��XO���A�Pq��x�����^u0#��*�g-!�Θ�QDoT������w��)����N�|� (=��v��XN��/b~����rօrE�`Ⱥ���M�Wq���ؔ����L��y Z0-y{��ng ��+��
z#`��#�����1{Y ��킠V?�a�:l9��@\��$�k\��kZ$�'Z%���٢�y`��ގ�<�B#|6޿Yx�'7��������y�ӆ��1��!yN��ۣ�a4&��T2X�#�_.�g�a����j�d�1ڵ�!M���3�y��@B����nt��ح���H�e�b���zn�V?XlxVHYEB    4284    1110�m?�u�݅�;��}?����O�	��H��ڌksX��~���(����dB�R|���3��0&Zm�jݚ<«�p�sLx��������5A��ݮ �>�A{���=^nl��`��Ֆ�V�rJ�Q]��1$#P$	#G���\����9�@U=�5��~�$�j�԰��"��+z�ʖ��?�
K��A��~ŭ�Ο*Ω�KR���1^��M�N�Φ��E�az~��Ek��.�w��k�P-n���?�먪�	�v��D	Ko�V"' �$�I���\ys�| :Zu��|;oK+;oYf�I��;�ӕk8�lB�b~n��
����;.X�%��g��'��M�ef�\���3=I����W�3
�:S�Q	Y~��|\J���"��=H�Eze#���8/᪢Y	�s`�\����G@����-Q鉞�l-��p^��4ڊ�iJ2nL�b �]=���o���c�1��Q}�ab"(����s����~��o���� x/���'w���'���"a6�����9��������1���)�:�Y_<�jҹ��cOq.,��G����Ѣ���{��G���<���JQ�8�x"c�m)��X���{���"t\���M�5�X����=��|JpB L��s~?K�M�e���-�|� %nB�-9���X�� �0۾J��#��V��g��!<�'	�xF�xl��� wS.�
Ϻ���Y��U/�G���D3���Qp��L��	X�9���5?�Rhvlf"�C+4�*��V||r���&��q�QF�75���9< �q�{ ,q9�j>�:�xԷ�i5�o4��8&>�,.�s��6K,�
��}�i������R��$�����Sz�L�6��W��s�Uu�R�~p�k���J2�|��K�\j�;��&|�!5��7���I!���G/�V�S=���P/��aV�ԯ�UQv����lH�W���I,h����/���%�(�:�wg��x7
��M��.0�Us�F�9�g�`��@X&-����$��	��=�1��Ā�CqJ�{�W�
�]ǆ ��g���b�⪟la�Zkă��g��HShx�+�7k6J�n�~%2C��9��t�.��3��F l�U����h�H����*�]ख��0O�_�D��Ie���-��ɫf�l�ܞ��.s��jZ�q5 �5��EE�1
�Y�p��61��Rf���$CS�n|�|���B��0��'��y4�Yo{2U���\��(�l/��~��;�Rp=�~g��@pJ�ᑶ��Go��C���/R��MF�-����R��V5�v2|��0�����c�2�v�ec���E����t�����2ўuy�D��
|�`t�Rnx��!�~�`�p=\�C.R��	;f���[ܡ-�I�$]5�<��C�b5�ٴ�%�[!���W�~�p�xc{�r/�H�X�^�h2�3C �o��|�i�杖A�[h.4Ct0-�_$;آ�7�I#|u�9s�]#ׅ&W�xKQCF�:��Q?
�B�O�覷8��0Iz��==|~t~�ན	O*�;�'��K��'�ba�ۊ@`�S�L���3^i�2�V�0�Ž���t�b�����|�^ I��`"oU;C|�P���8��k���^����i3��rM�A��.�?��/�j���6��C�xM�u���|�	��o���2�j�⣆ﺧn�bl;�� ��W��=��a�Uģ����}�D�P9}�}��8|��A�%^<��w$<7BŽq���w
�����B~K� ��4�w
�@F��L�]��j���{�R�҈�<��Cc�3�����{��GӜ�=*	�����$� s�H&�u9�R u�~�/Jy��!a6��9N�<�� =ʉh�o*��,��o�� 5�N��ˑ����1h�11�w��ړ6�	���]A��uFL���7�Sꗫ�Wf/x��nT�>��d���L<]��\s���*4\sʎ\���!9iw�����Z�c�4�L穣�K`�� ��@��z��3�v��"��`�9n��d�@"�E�Xd"-�@��l9����@��v{���wtP�	s�h �X|aÇ��8�`7�=���>�%���m�Do:�}P�͓�H�ګ����"݀׉V2�f�ʓi�u��7ݭ�B;8����Py'�_z_�
uQ��Z6�-W|��ç���)��꟯p�OJ 0Ġ$�GvcD&P�}��K2j�9v��G����Q�f�[�,-��؛�������n��JV�p��B�I8]L�I�c& �@z
���U7zצ0�X~Q�퉝帗�9��,�}zg� ��M�8�8�vm�le�?�8�k�*rZ��7�ѐ��>��E7!��F���>�\B��>���L��bK#E�W̱~���t�u�_v#O�U�\,A�:�_�R�g��)ۘ�K]�M���\J��A���HR{�HYO�U��yqZH��-~����\/9r2�<�!@�:,v�˸�3��uߌ�G	g�s�l���Mů�c�K��eȼ�W�vV������}'{�޷.<�+`.�<0��
�G�#hNf ?�}T����p�]7�y���D4tY^��`~P�Z[�4`�9�y;X���si�]�L�b@�P�����J�y��պ"0
���z<�Wė�A�K�����j�ʸ|}�[JQ�GRD��*�@Ѯ��/�]��4
)�ec�ъ�C���tR��J��/<G	l号+J��b�k�;��0�o3R�Up�b��&��QpS5�P�'?�t�
��R0!Nd���N�1����(f9�f�S�UV
�>kdET.����N�R�� wm����wX�����U����l0g���1���h�����2j��Ϩ�=͚�;��C0��^=���Qu��>tt QG&��)��t���IkYtVF3�R���Iy�3���z!��4�Z��P�P�p�Դg�n�!i�G�rTZ\�^D۱(�O���9K����Fҡ{BF�qT����\���з]�qC'��i,	r�a�v��[z�˓,�RYu"_��K��l��N���	�
��dQ]G�W�?���R̐�6�5I&�������3_+"��lT�L��L�F�7���6�v�@)�g}���C�jE��"
�P����&������	��.�?�#�m:���!ԧ�6�,aƤ�t�D����ȴ=c��%Ԃ��>UT���-�dj�q�4pg>U�0�Rf�~�U+�&��?�;D�sF���ݷE�m.c|=�������蚬�1[}�Mln")ר��(����I�ؚwt��Bu�����4H3F�!CHW���Y	�
n~>���,ޫp��=��f~S"�ְiޢ/r,��&h��̌Jr+��=�vK�cfpQ����"-XT�3�޴�@m+����a�E+P��RX*DD����%0m�x����}���vE�#�Cᢱ%Ϫ�&B���򇞬��<L"q�����)|���9kV�����`��3=�����k��RxT���I�]�����<-t/��B��5J�d[.v�,��HG�
۫@���Xn�V�TU���3�!��F�~4�;��N��ȿ@^���W�9*��@ui��J?�K"8����� �7�x��V"�Z(�����,�A��/Xw5� �6;��6&i�4V�?0SVM�Rm����p��2�wL9|ZPO��[ʺ��5�r��4e����A'ԝ%ΐ[r?؇�E����>! �zp1$�^�if��f�Qt"8U��=&�,*8K����QV�J�k�����g� �-b$7����ܺ�v���/ϔ3b!/��#�s�#�~����"t[)��#,Z����COI�5�Pѩm��A7�u��&d;);ܡV�AJ���*e+�C��< ����<�V��2�BX�t�:}�X�]�m:ОSh�y@�M���
�--:W�d�D�b1�>sgWm�~���*-�A���Tr�-�\?��vZ0ODTY�ݙw.3��'/��P�Z�Y�%}9������ω�`w)iΌ�Dt���.�=�S��̓2i9�[&k����7��Ѳ����S��Ix��zI�Y=9�
����z��H=�h����Eɭ��rzO�E�w ߖ�F�處֢|�?��@y��ɸ����H6p��?ns�*'������&�d�}���%�����=\	�t�������̆�WU:g�.�__z�϶��� sF�Sp��A
��}ɮ����a�٬��;�#���5s�PR��u_C
�״6xL�DY�g�Ǘ�Ƞ��zS@nאW*