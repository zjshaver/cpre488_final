XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��+���:�tv�h�:2�H@�y�(��D4�P	t
���w�'�Z��'r�8
�;�6�Ɍy�
�R�a�/;�Oֽ:��.?�)㞀Y[�ܓ���Y�}j�'/��Ӈ��i�W��r�P����QOÒ,^X�S���LL�f.��q�ؙ��ox��y4Y����� @�9*QD(o��n��w�S���o��MnU�XH4 !=�I~�,P�:t9%)�X^k��k��i�A�÷
;��ݳ���۷��*��9���Oԋ�޺Q�-v�T�h	�rppŢ��@T�A-�m������R���r��_M��VO�~�q�t�x�K��J�|/:N����+��z�ƴ7��)�Or���An���0��!U���%�!߸���=�FO5�5�@�^�!�}����L�}�i}�B��D���
պBu�O)͏���ˠ.���N�}���Ko�f�QW������C�5!7hI�j�\ҋ�h��z��ቢ��\M��A�=Ŧ��;�5�D��f�!'+���P÷�uj뤹S��~ -��ύ�񿰫�*AI����d9�wk���~%�Ϸ�s��\Ϳ$���1.�a{�3�ؑDW�PP�tcm���΋����f:e�k5�쭌���f��`��:b5n���Wn�&�d�W��c>�2��ə%�:gaJ�w +Č>��x*�	2�����w��	�n�!.��E&l��Q��B�UT<r���*���-�	$`r.��#�F-9�i�+XlxVHYEB    925c    1a60�m��Ix�M�F(7��$:��ĺ%�
C��t�TO���5�+x=z;�$_b�	�y��e��vAt�h�?--�د�1�Q�����q���KZ��i:��425i@�����7Z|�LP��5��8�(y��+�>�Ý*�>%P�Y��<�|�2���qP����! -�V������g��G,�]o����̀u,h3:��YQB�≔�GwUd�+g�q�z�7���;qֻޤ�N[���w�$�����c#�^T!�i��3A�
Xx�>���X�B�<!Ϧ�ۙ��^�WL���D����l����Jz��9���xUO��׵�a�Gl�~��1|�un2x�F04�`�����[��6��t$� �A�螶`�@���W��X�,l�{��2L�1����+^FQ��@Xs.�MF�
0�S��7JS;KNvN=g�h��zP�(Bz�)�)zE'�8$=?��iIh�LuE�dT�[���B?���Y���4�qf�Ii�7���Z�Ql�f��.��Xrq��v�%K�֎N��#C}�'������z�nda������X�y�����eO��n��|�ґ�RG2'O�Gϟ����b�Xn�J��E�Ҋ���^�$4�<�]<��r@��{L�=�]��@�(>uޡ��7��<f��k)8]� K������cI)h
o���jh��Yꫜ�><�Kn� ���]��v�@3�ݬ�,��q u��Æyөmt�'dE����#��7����+�?�ω���5;�9nCr$Q�2�Ͽx�.�r�>}N2�wȖ#&��:hc�M!��6JuSZ7%}/ͱ)�3_��a>�����q�L���\Cڝ��Y��Q�|�x��������]x�	�ݔ{����*>)Dm��0lߖ~���-H�w�6��޹5�C��	�5R�&��)��"�\X:��[m�,��ml���-��{1Rx]�5�K�Q�q>+�T��g��c�z��|�
e�$)�?�6?��%�*|��Bۤk����	�{|�z"ֻ1��I'-Z8�f���ɨ�I��R�1\�.�?K��0�qbR,�߱=8�m�u��Hə�SE�oD�m[탊;iEV��� I;H��#H)G���wL�m8{õXk�Aj����7�*�~]׀��*��?�t�2�̗/�tyZ%�I���*�؎�ZB��@�������>�ø�	�q�z�~,�������\[H�>{�r���ߥS̰)\a.f#��ī������F��ۗ��´Gb��g�t�ͳ��g���-�ҥN��m��L�v�7����y���B� i�Tg_��I��A�/�&�ҭ�^��9Z�
��hEg[L�������"C`��8�]�v��'E��Һ�'T�$2`�R�ǳy."�t��N���x������!�Z��d�ٽ�aވ������hy�asѭ<g�:)І�J(����Zc�m���BM��C����d��4u�V��V\��H
�2��N}���/mTG���H��C~���2�b��)6��a�M�
��H�NqO��A�4���^堰���{=��5������8
��%�~ZI9�Cj�Yڡxmv��נ�����
b��*0�������;��4�>r�p�d�@�A��]���j�C��w��{R>�`]����u��&�*�B��E+�'s����/{W�2�u�C�h����m��	�W$�e��p>��R������)c���Kt�:!�H��<�U�3z���_О6�v�(���9�1�4���%�,�BJ���比��kw�����H/D9�b�]��vB8�
��jok8�y?���F��i�m��5q���u70*�
�{4L��HKAvy��" ��'��wV���s"�(��;��Gj�5�5-3j?��3��\P�Z�M�*ƍ3Hp,vb|�F��W6Ho�'�I{v[�O�/O�lPR���/|�J3S�/Kk�lٽ���(<���xU�4����e<�ߟ=!q� K�U��C�*6,�g��a�����t|<#K8�Q�T��%w�1)	�Qj�`�챋VnX��X��4x�	��ݹ�)/i)娴<�I:�S*굋apX�`�\ké��]�K8ݚ�L]�ڐ����5������ܖ��%-2RQl�Vt�f�Ҷ��y'j�UW�	Ǐ�����niWz�����C�O���#$u�a�A����ELHG�)N���b�34��m�����H��-�-ǚ�8�7�TG�Zy��J��Y����|�{����<��0�&V[Od�6!;bp�|��P��g��W衬����� #�.��0`Ȍ�h��짉Ⓔ��t�9^�8�$؝���~w,��
�e؆�y��"]�szG��a��f��)&��-�O��yq�#��q���!�~�Tf��`����HWn,a�1$�˚��� �� "Vu��a���� �
��ڨ�nCZf����y�(����zn�8c_m��E9=�3R�T+�}����!V%D�&��Q]{�8��+�'�J:Iu��}�o�?��?&rغ}	Q��
�ƌU͵"K���'_I���êT���*зM�۶��m�*ֺ�i��vz�?ܗ���'NIB�����>z��*"şr�+�|0Ce'�%O�D7��'�U�V�Sʦ����ص�O�z�Vܚ�*��`�H�J���uJ>�Ƅ�}���:�l������N�Fn�*	��h���Y���l�;*�UYA7h}QT}L�Ƙ�&h��׾�U�p��+G��
���+��|�e�#6��8OL���ɥ������=54f����%97��j.�E��&����"^������I�����f�(�?���o6�)R�m^��8�	Լ�D��Ժ�P�RJ^��(5T��tc(����/ѭj�=T
1L�J0�=���'h<k��T�����c�*P��,*=��_�n�G���ћ����N�sK�{KxS��pw8������8FzL᮲�k�����6.*�n�	w�9���AWVέY�5�5�ST#�
�#۾�\��@�R[0�T���(�D)*��x=���H�g|ҋ��B���h��C���Z���4v` �9�^A�T�Xۢ�c�U�4�:hꝲ�<�����P�S*~�f}�C�BC��<����'I`��(�1��9�~��x'5`���e��T-m_�bȯ���q�S�;Gx��6�Fȭ�$�/��cڶQ�^Km�!�<[������9p"�j���D�ޖ���1��uşSU!���Ң"d� �����Y�+#t�Ϗ%m�*���ۍI�Z���1���P��݅< �F*9��A��W�H,䠪�,�i��a*'�U �L'.FHoI� =D�,:�1�X߇���ɤ��4�gve��2���%� !�����ޱj��m�AI搦+phD��߆�����될�O�{qq��s. �ڍ���@.1C������ �,;&�b���sDR'�(�٬��b�+DmK��6y��� +����<k�/��
U:�#��&�G��.�@[L��e]��<^�?�P��_�v�ߌ�ƥ�L�֛sv�y�y	���ؿ�O��B�n(Lz�	(j�g��w��{���
�Ir�V�)�w����'���S�_��,M-�B��9�@�gT���Ǝ\��A��:?W�<��p9��w��i��BR��[�u	;�˷4������j+Y���d�Ӡ�&��M��2|f�^�)KA2P~���=����_�ҢBC2�r��b�+�i?�]�9�1���x��1�&��/C&E�Rѓ�zX��#�ݯ-�5�z��!cReE*|[
)Q* ���	)3��yZ*�J��Aig�g�w�X�8�y�����]�:�`��f{Cʵ��&�4�;�q8�o��F(�y�'�J���<;��nڄT��@��h�v����K�Șh5_���E�ˌ)�p�� f�g+�*��e"�E%�8=�R%�A4�_N�L��#XdLFPLDL��b:��j��p y	���@/��6J �锟T�c̖���x���j�s���IyT�{�k*��\kbK���@��1��S�a��4=�!�	����=?1܍.���)�ر"����|�(a�!������|eL��K ���:zL�lX&3�my��� ���H]����+�PN?�,r\���((�=E|�,	��˯����M�g��z�aA_����>5	{���7٥V��@=R��FT�'o�,�,yv2�m&	&y9|S�|F~�猥��6h��H^1�tn���X1��о&��l狙����N˝���v"��2���t��	��g�s|6��e9V�{F������t�D�&�O�d+֣h�MF����d���)�Ӣ(7����
_�����j���Nn�l��O��p�B�߼���T���H��[$������0�ާK.���0t��$��YZѤ���|8 ̼p���C��+�(+_��9�2�����X�É��%$*^!s~�͍�AC�Yl��:��9l��ku�#5>��j�ٯ^i��-�����d�yxN�����D����V�J,+��<_�y�
��Pm����cov�L_ۑ�m@�(U>�O�j@�7bt�h\��B���(S���1�F�kؖ����;���܏�-��/4?t9�����S`QC`;��J��YY�S:��˄��n�z�dsw�%�GH��K�/��b2�k��K�Â�Łj�o���6;�D+������Y����O!�Q���E:T�J�������ׄ�2˨�aym!���ף�ү�C������,���a�Na��*��i#�Ӫ�[|k�𧴞�:뮖*�Q�L\�a9�m��<����P�<��e�P�A���f�IB|�MN�t̠���� �X�֭е0��m��9l+Vpa!,��)b��>�HJ��VnU�zbP��T�V+���Ȳ$Q��w'� BpxA�OC�t����6١� ��,E�(����E! w�h��׊��E��{ /@\=A����<<Q�+B�t��:���Zhr��N�c�� �[��s�2~�H���W�&�;ur����N�_�Ύ���ڨǍ�N��6�a{K
P�g:52c��	\�b�w������x
ψ�!�R�I��F	kǙ���e� -ݾٰc7�	�����<������6ɥ�F�p�����īy�S����N}48�}�#*����o�P��7:��%�uy�
���]%�i�� ��L��!:Ck���)�C㔖�bx�J�t��Z�)�?�������U��6 K�����u��B��ڳ�?�R����j�S�O:�4�j��o�,Y]�?t(��3R;�E���?������1��n���`Iyû!h���(��vq�����F�M�C����Nu��1��''$Ӭ��k�~�̂4F�ϖՇ|�"����HaAgW�ԭ���RX׮rIa�t�"�2�!iN�B��ԣK�s��½��������ő:�$�giE�G��)^�B�Å�1�I�!���L�|�͡�W~��%��H����t�����s�"A2�<uN��������o�,gT\���	�������r>��Ko��f��.�i���S���0����9\�t���ri��@�������ł=y��DHG�M�W/,[�2�3^����Y�re��[&@H�:d��lxz��2������QF�"[�%�X(��d�gU��F�F�wwP��*� v�zz�S�2�G�䀓By�K'��%�K����):*n&��X;u�q!*��=���l�Gu�K52��M��p��Ch�_����:�_ɣ�׳V�C%�	L�r��,DX�p*�]`a(����H��xNJ��J�5��s��'�V�i*�S����ɯ�����+��w��K�C�;H�fb�s��갶�T�HRp���K��W]����:M�}�TE����w�M�uڣ�Wd��%9u=���e��7��fE�[�58��}
��r���`��	p+�� ���a��aM���R�B���ɚz�}�S�&ϳ2�&������W�AN$��76Nu����.�3k���+�����.�B�����`��L�`���J���{k����D�;c�<?�Mr��Џ+��j4�v��m��YM�=�Ydn�E����!$�GW���sK9��D�W�Ց:��Z�)j��v~FBzw��2]��mVpߡ?zk��I_čG�)F]y��i��@}a��n�ļ���j������86-+�Dђ��DM>m�����>ۅC#OҞ��U/ˎ��?���Ֆ��e�E�Yn@B'EC��I y���%	u@8I��=1�Ɵ�6A�Zm[dz(��!�*E�����>�t�3[��v��!��A�����Y�f�V)�A�m�d6h6��3$��˴[-V!��]�
A3̍����	���3�����p�i^W>�nM��մ��ѳ�_�X��?���r?�k&?��\>Y?�k��"&ȳ�w��+�Y�C�g���������q#�C�+�P�e��8�>x(�n��+W��l	�3rDF���:[�Z_䍮R]���&��I�λ� �4ce:
T@y�6�z�o%���|�m��b*˺��i��