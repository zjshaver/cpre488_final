XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��-�6�0��(H��t����̎%3#a27h�q�t���u�c-Vg�(�w#@٨D8S����Kqy! VK*6��qx���Rxľ��V�Q� ƽj+���1��������1�ܚu�2Ԕ�w��Χ��cvV_��A�Z�f{Eh��HV��G� ��v�\ڸ����X$1g�\u�5*��C�f��1L�v�sb�oVԴű�ʮ�X���jU�X��90�Q�=?��F��,]����_c���ot��I,�Bh����J�\������(�v��]�$Ą����΢��IW�|�YHu�1y��9����[Cv�5�\���X�8��G_��l���d�`� $����(�����wg��yLh��Ak�w��Uo7�������DbP�� ��[,��Q����fƐ@^5�z���/�0ҍ�:[˺�H~���)���^�B�yh�|e'rT|�_s����|�`9���x�nU"����tk���,�3���	g7�a�>ŏMF2�2�����u�.��N�����"�oL=�`u�B�9W@��$~���w���IL�5u�j2�1�Vp��zQ��� W����f�p(=h�mV�C�Mc�O�q5�� æĉv����^�X):�#1WU��\<�Od�e�Z���c�zȘͼ)�j��6�X��d��]т~�QZ����6ź��+��#r���'�������H�7w��tё�hcx�*g���Ue�D:�ǯ�dx2�]��'ə=)B�i��r��k����k�27|XlxVHYEB    7265    1660?:��D��R�z��gLT�j��a�~:���N��C�?&�lY�X9��a���E��nΔ�	2�1b�#��9���MO_�@v�1�*9�F��[=�w?�?`y�X�m�3��
���+�{ܚ����u�_sK|�L�5��8���;��ɢST͵J*�$ENN�f���>0<Tw�K^h~6�r:�6�c�@7�	� ��*È5^�+60��3<�Pc�6�M#�ug��b�����<������S���l(�? ڑ!:K���A1�[cܝg�����ҩ&�u�*����ަ+"	�~n���@�i6\��j�<L�*�]M�����iTJ]�i(AD��!�g�\ѧ�`w��LJ��
�H]�IV���Q���=�P٤�$�I1����r�-��o_y#�p����LLY�#��$�_��J��?F�������ˌ��=^�^~TU��]�V�:�ܴ���5L��r^�@9�������6w����8���oMѡF����t^İ��`M-W��F�� b�]ˣ/}����R�'yL0d�R�/�C������!m �2�A�Q1�+�`о�2V!�_��C��YY�&���k�}N�ϖ�������_�^�8��qZ%{�n'�v��A�,�������*U����s]���Q#�e'���5�k�+v?�;"H�6,\QGPHu�����7� �
~�i�c������R�b(��9�d�K�O*(|���bX�ଏY~� ���a�$Z��g��UCޛګ#V;�c��5�z6H��al7����ͷ��U�% 8�Ux�<p$��������u$���Sd`7NAN��� ��t�$M�G$lw�
�!���<�������8���@�&��4��^�tS]m�U'��ͦ��+�!��\�{�HX�g7&��f���WUC��]�W㓞���o��K1�y��M^���&;Ǖ��Ւ9�^Z�Y�r����P���k5a�7&��r����P���]�|������lJ�)nx�,�|{G��x��0Ph�P���uR�!1j�!ؑ���EZ��~�G�b��gyq.[�yCЄj�0�_	�G��?[�J�]T����H�MH��v<�@(�0�A�	�g#l�N
�ԛ�/��26Z�VK)�~i��5���B����5�rJ]�R��*����wDU��@$ |8$
��kB�����u]oFs�V%�M�_��q������H]���4�_Q]�Q��w�u�sd�Z�� �%8�N��B_�����,��j�甮&J���j�J�8�j�U�Ug�.����{��!8Q���D���R	sD���_n�^�	����W�R����ĚWb�����ݛ_��P�X�%���̔-}�-���&`�	����h��g�f$�.<N�>G�~�����4�\R���6r�-��I���O8'���K�*�߄K��eKʃ��-5N��*#���[�^��.��;�lV��nT���i*q*�\���%m;�2�W勤 ��	x6��Y>#�h��G9̳��몫��^���D,t��:gmt�2[2��MR���|{�/I����υ��!}b��Uw�:xv�}��֐�#.��Jɡ�=��7|L�	�o�1o�$���\������kfb2�B��oH�D������'�ߟ(���m�X!���K�����+�����5ҍ8�VTb:sb�Q����f�"V���E0O��~�Lb��i�+�/�l��/E:���SWo�	��r�Y-��D�9���o��$�X�x@��M��s(=�%C��jo�k�,�F�$kq@�kW2��A�S@} ǐ��8���*��-�o:�ژOf�ucrf0/�}�#φ��x3���ܭ`"3k,7)�.,_�m�,_@L���>J	:n8-������3P�d�({�X���ep��RA���i��f�e�q2Tfy��,l��rr��[��]Dq��;���+�2%#l��}�ʱpC���!^濆���y�U��D���Fw��>m{�K�QuSj�^������]��2eF	�h�;3]�ފ��7�߻��$h�	iՐ�����@�i�^�#��t����L��w��ѭI�,Ze�|�儲��MD#惀�c_���5]�f���}ņ8*�ɰ�w�d!/�~��c�Ḻ�K#ܱ�NN_ʚ�ٟ�G�a�y��0�O<�X�n��י.N��2�oP��sOV�����8�����ڰЏ��4=5D����_����c0Z����tgm"�r�جu�%׍�t�����Yu��G9�cxb�	~�G�S.t��c���C��?-�@�l�{�(�be����կ�~�T�ؐD��%N3��C):I�aE�? Y�.�RˀN������W���<����� 5��`HF������@a̩�G�����u�z8+�@�Ы��������8,(�K�I�ƙX�HDK�b82�M�6��|�i���PU%D��mS�J�YmB��%H)-a�'
�z�?u�Ϫ��5��1��d�#�T!č�]����M��Sðe��w�;9�B������p�G]G�QY��4#�bQ�Սx�d���L�����e����|:�4������� E���o��?Y^)��ۚg�
X������HQ�m��R��m��W_j�ӆI#Q�(�oSˎ��YQ��}���7Fk/v���~�A7��x�: a�C��.3H���`0따�3���Z���^�_0����SSVq����˧''H¯Xs�}�Նmd;��7�]L��)[���-������M�ɉ��.�6��R&���;�f[@L�'D�l�8�tc�j0����� 4!�l6��7�$ؖ�
S�.���?��6�Qk�DV�s.mz�2����G?� �ܨM��k�tV�v�6�sms�$��HC��GQ�%N���Z�.�zKl��ɇ§��"�TF@*�>��釾�Ch�7�ϓ��7��#���b.�&��i����PÊ��k択td�3g
���f4�}���L{t."zsp��S�(��1b�G�37���;��3H�mk���%MaH���7�$�p�����4ϣ�(Y{t�=I�}�8��@4jtJNMA+�}�w�*�Fy�f/�L\�&a�#R+�P��g*Mx���$���?��؝��(�Ex��[	�R�h���Y�l;�E4qY��Q�����Xu�QcOm��Hgmlۊf�Y{�H?�6�aU��c�Nj$�/��~79�ã���	ܝ�@�D�u�7(�'պ��h�;Ѽ�sMpdĆѐ������4�$��;�&3`?6�ӗyJ!���c����.�¢p;��^�_�,��$�ǅk��t�8CG��@4�'��Υ� �6�gɡ\0)����0<���e��=��vh���Z�$H�$��PY3E�� �϶��>2�<(�n�_�u�V��^x�������*���-���&�밋�Y�p�+1��Ua����R���Kׁ�9�\�ףA�Z���p�<hS#.��l���i&��W�mi�U�5�ȩOb�X�����'�ޛ2�(mGf��:@�<û?T ���M�A�gP��\�b.6�gtO�{'��g�Y�&��ↁqC]�Z�̘��X�w�9�"T)5�4n/��5�輅Q�zG�?zûc�� ȍ$<�9Á����p*t����X0<@����z���E���[|�$������ʓ��vO��6��zr�����(�%��A^��8�֗�]�y2��t�mry9r�0��ªjX�$YBS��i0\�^�2S�
��
x@.(7U�-�>�L�8V�fq4ޭ�].&�fv!��GC{��f�q�f0�!�F�A����"��4�V�p`%��G�06��B{�;(�|\7"����{�m�<��a�Pg���iτ�����]ɳ��Լ/p1�:�'��F��� oH��+p5@��雏�$5G�[���u�����鍪���xX�=���܎*��|���~x=�r�
UF�Qז��D�����0)�ۼ�� �jz���f$���'�v��~�N�ٮ���Af%L��׍�`ST�?hѧ��k�up�wS@W|� �����2!ڔ؅�V�tQ��0]g��d�O�h�?
���� �N�>�H�á��t�a?&�Ap�N�6o�/���%ô�H]YB��O���1��]E�p��=e���%(m������K�����{���2��*°�������z��������t�m�����p��%y63-ى� B�������9H�-MY�r/�M_��= }.�w�;qa�t��C֋�aS��m
Nm
>~�S*M���l�G������Wr��O9rMz@���	���/�c��m���_f�'���gU� ��:[�c:���+컾��J�B��ӿ���?�Ӭq�)&�0��q��&amI
�b�=_XR�m�]���44[�����C�S,-��\e�Y�-��L?6�o��R3p��}�'�_���\,���N1��a���+��}��㚇!�M�Z�'�V��8����s~�i߶G����0 <@�K���y��eH��Z���I�����?��S����
�)#����ZyQ��@v�c�ي�ǁ� ��x�!ʹf�u��0�k�,-�Y�H�w�b;s��\���h��^������#>)�r�I:�f�/	�q�����%%�G��
��_����.)�έ�e�Qb��x<���&&ZV�|qJ��y��m��޴���@0�MI+ �|v�H��jm�m���}�R�����ϑ�/���{�5C�>]�	Uo5�fa��2A���1� ���������6+]��c��<�#��C��v;ƨ0N�̎a�g�4^c�`��O�{���}�}�| &���[���/Ɗ����$�Z�pGT-�xh��q+��;��n .��3��A֟���;Z2>%�k���*FnSK�FQ�������)܏�i"T_�������/UD�#����RH����v���I����5M�Ƌ׶8Ͷ����I�I���n���nP�K�Нp��ݥm�P���Է�R�$��j�G�L�'V�W�Z�7��*pƧIk5�&��U��f�ȃM���ƹ[\��k��L�!�v�w������o�λɠh�C��U��=Jhue ��"�U,�E�%�pl,΅�E��V������k���Qr޼���Ԡ��j0�e��:խ�r��{*�?����\/�0,ޕ��X�&�Sх!�&�v�����`8b��*e�#\��lQp����;1�]�A:@�0�OA���}>��(EC#�N>d��c�a}6t�]u�op@�W9d�f08(�S)��L�����6a$�Cw��_��F�����n7�%à�z����S���M�Y�8D��N������� $L}�rHg{����t�_׵N`{)���ڻ�=u�4�[�&7j�"oX�ܓ�ؼj���}��5����r��2p$�����bQa�"l�Lm�=��^o��M~$�Gd!Bր��Bj��]C�#(,�ۣcy�!93fx_�P��+�W��W��H�J.e��چ܄�3z���t��<Cx�UiǴ���z޸e