XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��V��p�\_���E��@�ݍ��NTO)��(t���D��JS�2NHD��q�6��E�-F/溴v	��g{���2�y�kQ�n.�Ae����H���{FK�?c}`�B�+�Ю�1�R����i��-M��Jg�r���[�Zw������l�"�F���7L|�������З ��fڷ�H� �Π��'�mI~�#�7��FB�}D�df�z�f�^���e����� V����m"Ob#Ҏ:�g~�omNt7�+3�@�ͫs�2����`Zk[D%s�OW.sn(çh�[t
�э��[�,S�ΏUY܂�c��GZ�k���\��E��&6��5�ys��7��wچ�E?PE��2��Ah��y��ߵKf���s�>����P"�^�ލZ�.	�����1��L5J�I��;��_��k��:�)TH`F�X���hW&,L#�:��l�	|x�]�;޵��Tڊ���zl�/����$�au!�������쿝����v�sF�&���4��f�R萒�p��A	�X2̪Y��ēTK���ɌkgA�8%��Jg��������I��p���iI�`�F�{�g���\�*E�S�p�S�NƗD;���e�t�Z�-�+�͎���}7�}�'&!ܮ�'��Ă�(�6#O��#��m��=��x��k�Eo����C<�ƞ�؃u�oǰ����`Ix63I�r{�^����n�w�����5��24�����υe��Hr��/�GƟ������q�T�Ӟ��\)��XlxVHYEB    1959     920�L��A�16�pOE��#���?*��� 5�?��.2iv�rC-"��1�7���a�9C��g�LЋ��)q���)/8{�&�ÄKy�*��*��"���'��O���y��� v����Q���e� ˝�
���ms�u&x���! �&,��k��ǈ��|�%�<�e�	>ZѻYj�d�� GKw��m'+;ۑ���(��4�ۂた����z��Z��m��B��$t�
j��ǀǲ�&dk}	?]�, V�͕�]�h��־��?~�6���M=_��
�a�ډ��#� �M\έ�.��`��wUQ`{f�V���g����`=[���{;ߞHP�e�|��f�-�9�֜%��Ͱ5�$�g�f�/��Â���ж��T��#��tX䅺	}ϟO{���I��(0)m�����`b��À��j"5V<����DA�N�a�	\&p����=��W+�r�?l�U=�fˍ$�g��V��hU"S"`��.]/�fuN���~���~2���T���SD8��Sp��0���л�,��۟êwA~�Rĥ��^i,��V$�n0}I����H�3em��ҨnϘ���ٓ�2Ydg�x�	)2Kk�B��}�0���.��2q�� +���,�_��@����Ug;���VM�����(J��T���=<]6��\*�������7�a���'�'4�!�|�+Png�˳қ����iN����)�x��0�TȜ����=a�M�6���
�6�����Z�$����(�71�POGd)� qB0<��7�0�H�����?̍^��|C��������j���AV�y;}G�@L�s?0���l.X�)�)�B�ڌu��jӇCD3X���.���Ș��inN��l~���B�J�g���w�����[�-����)%���Y���=6B̙+�\Yq�'�{buT/dy�=e��^%^'.�Rwv���1�b3𘒘a �S�˨:�ٟ8jMm� � 6���0Đ�y�Gv�B\��N���K�dN�D=ܛ�3*rn)�q��yv�m�'
 rD5���zs�����TB����N:H��R����4/!��w&�(�e ԫ�stҜ{l�7~?No�hE�%�N�X�h8Ju\	�t	��)�6���(�ɇ����F���B����a�E =����U43,�G��g)�"tv^,$O�%��W�iǽ�䀱:�'��h܁tg��D�f߯Vj����gd!�bb%�9�3�i��Ά&�Wd��L�5�(��c:�8n�-&��4PC�<]�?��L݅5�����=9U>E��xh���;���%6�=C����Zn� uƵ�~��2Ah6G�ʗ��@=h��ů�c}��.�u�mǹv����?v٫a��P(B��s?P�H�p���U�S�W Vuc��"�IM�,���mɌ���-B�e���q�w9f�.V>���Z�p�GAQ�)�y�o��sn#����#���^�M��|3�}ͬa���Z�.���@5l;��|����2���L)��~0�9z%���o���]{�[�>�o�\�|�M9S}lu��B�D
�%��vs�J�.e��j�����٬�Y��Z�LE��&i@���0��N��@�[�ʧx��;�_/9I�p<K,A���l�m����T;��ձhr~h_0�����y�$U9-��r�_]d��KJ\r��t�a�	����~���v_)f�B=����g4txDq��0�����/��2��k*�b�HeK1��/X�d�v�LTx��jњ�p|�_ɳS^	�f�+�"fe�D�:�Oa���ޖ!A(W�@�l~�a�9N_�.c�	{m8tld�����0�q����2G(�*��U�֌̫�9���믢�C;�����Ho��H����AZk�9��1C��Omލ��lM>����E���`�7����n����}��-DoN��Gl >���g�&�G�b&E�}���=�SYh#��w��Bn���� 04�}b�?[�8�����oT�@iK�����͐v���2�K�2Q�\�7i�Aϋ[�;o�7��Xx��n%��ug5{��L��u�Q��̋<������eC������:���竍˙�^A��|�#�Lk�������p��zKJ�vN#\���� ���v���s!cf"��T�'�� &�W01@�$!񀧍��7*�w�|�V���Ҍ�ʆR.��?h	@._$���j�W:�:ß)�W/�#��ab�Z)���}��G��������>O��!�O�K`�(����D�