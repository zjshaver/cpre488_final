XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��+Jn_�	���T�����"�䟹��)Vp+Ty�O=Qi�������3�PMlDHqƖ�䶻s0)���5�vF�th:��o)�����j���o^�~�J�8��1=�ӓ�J	mNuB�#����O �@�p�͜ex�қ�t��rI� u���B��C���~D�?����"���$�'����>���6K3F�i>z}L��P���T������B=�$��9g`2���b�s�~�� fDR>�щ
H�A��ڠ#�p�:x&�V�D��O������\�{$7��uJ�U�ːKܩ���P	�?_�&=�1S���W3�(!�G��Q5�Bߚ�mQBL�ma���f�#Hx�[j���ӓ��-k�L}�.[Z�����~���my�շ}pv�O�L̉^�x5��aU����2���X ��+�g�a-�N�������A(���z;���;����!��~A�vv�?G p�v+I���5��w.���fH�1lά�7JA�tN�iXv���q��ٸ����j�|r����E����m�O�`��w�,��s��w�WC����� S����6a���J�[k�J����.[g�C#�"#黷1���1Ɖ�04�j��k�<I25�/���*�F�\���\�c�d��	�^��~:x�FA���qK�t�W~�/R=�yk����	x�"/�
1C|>Q��^�m6ņ��N�8��ǒ�_�ڃ��g71���};XnR]�����幑�E����<�ZGOXlxVHYEB    1a2e     8b0�j�D��z�e���+�[ �R��[�����MkJ���A~
$�}�J���T��fR�:5�5j?�����Hsb�=V̳_^� '���|F��q�b��1h��Y�Ƞi�gw���ի>v�L_�Ӽ�tt��>�ae��Z ��# :�0���6�$6]n���rh��%����`~:�l��� �4S�j�|�"�Sj��h+�7b�5��š�q6Y�P��B��\�<40F����nE��Z��#k[��X���H�+J������a1�6�����/��Q�b�X�#v"�����3w�u�qj�c���p���%�i?�%
Au�n�+̻�U1#�����г'���@��'�� Ox�t%j( Yn*���y<_���W�0HYk�;��:�0��*Ϡ�}Zj���Ɔm�}�dx6s�S[6��͡o�CG`v��z�L�o��Q�O�3w�v=Rs�JR�S�4FΤ�Y�v��/+�P���~��#�Q��kUQ����V�ƨH���s����:���˓�~ኹ����=l�5��N����0ɴ6��ʃ��BC���$��X]�m~���hK�v����o �7�9���/�R��d��GCͶ��:nO
֯J���M��8�ۂ-��l`��F��u������h��  ���l�ɭ��PkE-�R�w���3�m"�i�ܮ�d!on%l6�ھ\s+���홅mـw��o�8���Cʣ�s~��2A�b���֓��+ϲ�"�(SR�>,����P�R%F���q$���1���2>�����T�����E���&�탒�����-2�6��eR��ߧ5��s�@�YO#<����B���_Z�>�#a+�8���� ��}Xܻ�ĉ*F}� �RS%��ON�D@�F�}V������s�Ѧ~MZS���\.}1Ԛ��p�D��/c�ܦX�;�#&G�GN��������Fm]cNbA�aî����8~u�����k�m����
A_e����_l˜^q��Y���<ɝ?^��M;��4Dt�p���Ƌ,I;A�`�v�%񒼷%v�V� Z�`Tؓ
#�5|q�Wn@9y��,0��#38_%# ��9���B\��o�s�m�(�x��ly�;+.���H�`ޭ����y�p���н����X�
OKU{�;��i�Fb������ ���
��Q�n���+��z@tD]���V8��n� ��dR=��b�;�`���*�}�_;ۆ�[>��X����$�������$�)��Y[^,�vU��$�XzP��'���%a�Ќ�몉�� Ώ.����N	�L����|��B�J�	���u��u��Ϧ���WP��ߞ�w5_\� [����30�o2�[�Ω ��R.���*��jP'U�s�ׇ̽��;�A�GZ铸"�Q9|1%�L�"�ѯ�ś�&"A���8����O��J8��!t�5��7��f�D2W������Ҽ��+2cx$?���R��C���.��$��h�&�8��~T^��Ѩ�a��9 ��������g�|iw��"oB胰�f%܍)h�0��0bY�fl.�������PQ9Oo�]�������#���&#�����"sl�ð��_x��0j����~�)9֜�)v��=Ֆ���⃱v�υ��X��DC��#)����>rfl)?E�e�׽���%=��X�^�Ƚ�_��uS�Mud<P	��-��Ȏ�'Z4�78���+��_a�}�X�����pt�|۵����)�l.��~�躭ҏ�E��L��.q�D*Mۓ��KfDAb�S��怾��]͔d�ݳ��>=���e[�u۹%�r-ⴶ0ߛ�{;w���7'���aɷ�>~����Y^ጛ��3WY:�F|��>��|�Z��ل<���U�HmbV����P6��,�g
�k��a����0�y�����i���4XҤz��݆�L��V¹w���3�����=6���-�|�EbW!Y6=����V��S�Jhc��5�+3�-�1�Ȟ�_=��r�[���ܖ�{�%Z�c��q�8Z��@�����J��k�L�׷�9 K�w�#�V��(N�%���.�Aڠ���X
&��=O;��<��]Má'h���;<㙆��`���软�4~L�Á��tF`CD���'�!H�?�kv�6y��R��y��wv+�