XlxV64EB    39dd    1170����rv�v/�p�u
h�Vf�`v"�r�Ha���m��#8�=�M��	r��x����*I/[�!'G��2z ���WT�������h^��i<�2��6����=n��8�`�#ȹgQ@G�Y
���)4�-����:�y�0����X���}fC%.��dI ��4C�nZ"i@�h��uT��1�G�nD�m2�ވ�$	�'n�`?g��"�������g���GK[&8����r��	���<h������h�ɬL5BN��և�M�r:Q@dxfY��Ƶ2F���d7�r�Q�8Q�o�P撌"��d`��!�I��hǻ�d�[9rO��H^�:�f��_$�"<dn��Mҧ�R܌ց��n���h��(q#赀`��3s��_H�y�Xh}-��BkU�vRJ��~����a�5�Y�/!��t���ȇL�	�� �3sp�H�m�0A��ߐ�{�$��ΐ�_IM�ľ�刉S(|�����/1�v��f�
F��	O�N��f��yEw{=aNN&��^LB@2�+�F-%�c]z�5V�����2r��������Z0ײ�.���c��� _ۗG�g��l��1p>��#��	�#l���ZݚI�Ʋ�����hZx�$6E\��a��g�[@�z�/��{��u\�L}V���<C&���ٔv{W�ƼE t����ʀH)���zK`�o�y�2�H}�щ������(�]�gIaw��$'���XjB��_��;��kȦ�O��0�^X��E%Ӱ�k��>���k��Vc�B������zu3r#�H]2�nQ�Ǔ�=k�B���Y�T4Y�U�F��N9��0����;��nIS7��2垂ꉬ`����g��Ξ4Y��h��i��$�ZN��C,�x}�:D�T52ګG�s�/���M����Q4���U���B�I�_��}�C���
�΂��1{G�̡:(+]�g�V4�V�(l�DBf�	�ƿd�Ȏ�m[!�5ãhV)]�OD�I������gz:%���MOs���)w䥗!q�Λc�ы�B$b�1�k���Ex��V��$$4�Ǥ�>$�[e
B�Zk ���� :@Z�f���O뫬��?���u�D
j�xgb�E�<f�J>����+`��b[�p>���%����;��[ �)��j���k�
2�y� }��"���5q�v@�L�g�}�=� y�����ֳۨ]���s���˺�C`��6y���RhU���G�5&�̜UN<m�����(L�Vnw�yݿm98n�<��'�"mOC��J�|�2Xbc��7�F�d�=b�f'Rr�Sr��bO�.F�vD��t7���mۥ��y��������z^m�ʰ�y21Wq��'"�ٯ8e���#(�GV�\�#.��R��"?|�|�N珇о� yQ����A��ʰ�M��}g�1L�X�6j�Q���\M�a���CCL3��@LXM�b��A�,c����(�>\С ��CU[>����#Y_[@���1�~�8�Q	��!
����5И<?�^ L=M/g��&��Qz]9�̱p�u�1�Y���<+�2p9d+��f��c��q0XRr���1�=v �q�:���.����c4���!��x^Z�ƚ�*y����aSM�+��͟��V/&�c5��z���K��G�dH�ܽ�?lHU|�%�|5s�q������p�ū�'K	q���Ė����%|L`AS�8y�JYs����uj(��{z	e��\����DLC	;��,��(���,���_1P���8¡��"��RQ����"��c�Γ���r~+'�����fↅCIK�����m�o"��!�u�#��N���'�����8"=z�t��gs^�]� ��ǀg���L�>c�R�Ka�&�̈͊
,Fޑ�<�ǒ���ha�_�iNc���f��p�/��ڑ�w�e���	5>�;����Ρ��\}�63��uj=�W:}�>���==I!B�40��I5�O��$�J���Xp��!��]b@,(��I[3�;lֻ9����[���7��cԸ�M�&y�%��p�HD�����v��D�Y�ע�!
�9�(�Ǟ#]���G�+o�T�E"�W���-8c*3%|�x��?-���� f�6�x�t�J�񅪼3'������m�&�&e��#��귑�����0�oh���G{�B�CNM��_�u���G��ђ�Q(���R{��j�_��`�
�U�&6`<�)�K�}z鸤�ؼ����j��{��Bs)�<�y��N?��]��ۜ1�#k�����|��4����u�:�*LC�ˈ�2{�lM�zA��&��H���س��O��xɷ7
�=�G��C��cO�;�/��i
߅�XT�WҚ%X�L��o����G�1��dIJ�̛RZįI����3$g��(��IN3Y����M&z�^˭�p˥������2p��.a̓���5�v�U�d�=F?V���;2L��@GW��&4˯ 3��F7�T��w��,��sԻ�]º��P9_��c+�
ܒ���nx�[L�O��@r�'��/���FN��鞴v0Rf�N��ח,����wODIߧ�θ*oN��2+�\�*�3�x�#.�z�}��]MH4pR���OD��)���.|�k��-δ��ا�e�N�wC�[���q���CgM��M��W��1k�b�nv&�k�*�.�@��)�@^�p}K>��O��8��J�ǁ��
�,���ͧD�~+a3O�p>�d�#�����st�����^܆3jX�E���;ꙉ�,k��
;v�9�jNi�H�
�,H^U��&��ż�W�kA�-c��<@���&�q*c�!د�h M;��z�ղD��/�D.x"Kz|6_��W˔�A)v���L�1,d�MX���a�XL���b�<W��pJ��J�-v�y��5Q��)�{.�IRR��k�
SnU9'�¶Iq�uNu���N<�6̲�bz��{?�=�bR%k�P�31�ٮ�3�����9{�a�hR��:��`���&�l
��	��ǹN����,|3'���Q�z:�Q3h�J�|�r$���^,
F��fn�+��5�>u����2S���r�H���P��K�а�B���a�o�մ���S���uW&P��Uu]�G�ߌ���(*޴�\�oF��V��;�����sl����h�15��i�G��a�!Y�\����.��DҺ��������a
���r3D�B񫪺7���;�$�u�l��D��}L�U�jc�һ�[�ZxU7���ŲvA��a��5!�_���T9���W���`�[b�\n���VĜ��&�©d�iu�M�FT"�wـ���k�/9�:�z��ó��t}neh�5����H+Z!>�<'���/!� ��ϵ�3V���������~\��7�,���Ī������x�Ӿ��[v�d�\�	���P����Ud8S�ak��x��,��d���7'x��z���Tyk�Q�:��w
~Uϫ������4�i�Q���6M���%o�#��.H���H��K�w��{%��e�W0H��@���������?���n�p�\�������$p�4����o3x�п{'�zixR������)>&� ���h*7F�?Y=�3�ᙃ� ��I8q.�!����
k���ɲܕ�$U.���1�T�HCN�w���͞s\�m���&��KY"�"�0�&Q�Gű��ţ�����	�N��WL!N^0��1�n�/���~�a#/Τa���5�� �Or��7B�������|o�P�����"��4����VCv�����[�x]G�gB(��>��l�$��4B��,Fl�;�g�_u��B���+~x?�kF�Y*ٛ>7�g�ݴ�lT�):�ƸF���xJ@uϔ�N%�:BǛӜ����Ź�d�p/�:���yo>=�M�s|�o/��ᖗ{�|dɻ���v����Kg�N��?����A�V���/i�'%�>'�,�榽o6������2�R�NG��b�(4�j#�DA-v�qil;���f�Bx	2$Y��3'
MGWs�A�d��:"@���{��g���i(.�h��Zc���;�nY�5Paݡf@5-��iFd���f�����$����.�벃���12\��(�w��鱊JR�}~X��J ��
�flX�p�U�~��}�jv�b�彺:8�ڨ�c�Th����0�!722�/���e�т8w�H�u�>��,��g�t�I0�i�
J3����*��"ڦ;��`y���_v���ʆ>��\�ݼ�v�c�5qewJw�ٛ�����Y�㥀C��n��lՋ�mh�86|��0�ו��2/��