XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��g�k�++ hgFJ5�������έ%��x	&�J�jP���J'�O��?�6@�� �f��i�/AX�vkUͱ��׶�c�dG�fL'�qV��Z��l�n0����O�T�p�e���� ��U����9$K�)���Ơ�:��.'@XhNxqS-��xJd�8: �P8_��� #��1*��BƜ�5��L�s�*��Ik^�)��8���t4o���� �l��O+㢗	f"q���V�|]t�uƹ��|������Q�l�5��U]�8����6CKB�P�!rn=�聛�'66�c��ׂ�4t~��_T�6*��
��9b4f��Ėw�i�C����-_�z��'։��$n������Q��0!cb�f���'.'NA�m���&>l�	��_��fYO�������eN@���� ^���Xףi~�1��"/"�G~p���,DO��S�7�Yۍ.��M�:;��=�ߐc��nO4����)l����ك Kv(DO����Y���� Yx�����e�n��C�^;M5�[U
&�5MyApB�H'���YW��V����^�������Z�Ț̐��ڹ��R�Q"�ЀQ�ܗs�Na�۳I̞�����4�c����q/��%���TB; �C�1(ɰ�et���q9C�=NIR	�	k�8���\0u�u�x�?����Ib��"
Z���$9�G�X�S
�p+?�	;H�Qd��a�W����� n�G�Y��7czv` 5�Qފ
]#4"�2�TmXlxVHYEB    48e3     e00�Z�S[�.y�u���u�'*�@�إ�`��2��V�ҦA5L�����5�Sy�a8߯����/=�ρ Z&�3�N�����ȁ����A�@�Ը����z-��gU�� ?��w''$���� ��4�_\3 �Q�r�3�%YԾ�����k.x�,���ó�v�0a<`��p�j[�ɿ��G�}�ܝ:�a�p@�{U,tRSr|q}��,���|�9q�B�E���Ս�Om}��`����m#�$/��ᐉ46H����ca�̮_x�@�:�?�/%"1uA���0s���ز���|��d�����Y�jZ�6�.ń6��Ћ�;iR	5��r�.����^�<��������R���AƋ����
�~j�{��Ix�����#�H��z���:>� �?C�v�TF>���l`��d��ٻ�^64[=5T"�+D�g��l�t�B���2�a��#��.HZ�����{lF��o�0�XXj��x"|���"C�z��y�h+�:�b��e��}��U�W'mSo�Ō�lz�5ɭ��ڬ���ڇi�%�B�:�Q���}�_k�!�%��2����ֵ�7��H��#�F�f1a������~c���W�-":{\�=
�[�,<�!C�bp�w2��g;ч,��� �/p<��$ڪ���U�������lj%�jk�H�"n�(�$FQ�~>��6���v0�'�q5�Z��ϵ�T��H��� <��2j,&��c�O;���x2o*�U�td^s�&<'�{uuĳ���� �I��b�����<q��( L �D�4`�Z���ӏ=�?�.x��0�m���J2Da>��W�&@Ր^hy���N�o�eF��=�ls;��x$��a:˂8�u�&��\9�vQ��$ ����?op��BĤ���5�s��h�+���uYs�j�7�}�sL�cI�UO��7���U�Y9����:K�}<�g`����T����&P�f����
�*V��V�}�0ܼ��~Y��ޓ��/r���!�+V�Q���Tɶ��N��x�~�u�o�qu&@B	.6�NC�f���S0/���.��$U�ɣ&�-��>��q�s�ӵM�$�����B��G�oզ���woE��l���AԎ��	B��M���M8FM��3����#@l�x��r�m�_��@�ʖD��]�#�:�$����߄1���-��j\=A�x;CG j�9�`���8��`�\� .f^�#)�&��n�-	S����+׭�Tʶ�Ls���L�Ԕ�.���aaP{J�:
��%#Y/S�E�8Z梍�n���0����b���]�%����:�{�����qВdNĠ@�k��RcG�C��B�8�q�{�ud�d�10�l�r�.�����4[��w5?.�i�ʩ�0��**~v�8��P�cd���4��6��|&-l����� q�_9���������lC�(����̖���jaݠq��!����r|3x&�Cm�ل�V��)m��Q���fV&�E��k�s��6��<6��L"�����b�n����`��3��h� TL�nX�=���Ѷ#�E�hf䰏�3�G�u��hD�х��̾�V�4�+ܼ����@Bh{���j��Ħ��@�-��u>���t)5h�����膵ީO�'�攙v:��8�%��}���$)f�^��3�Z	��ŤK�-���y��z�/�3 \�
��pEX݁��~-YTs{�4���o���B:��N���-�����x_ʮ���=�\��Q I�V�b޽ܷ�^�5��ٜDk ������׶I�/�9%��0M�5�zH�h3��(���uUU��{����|%�tO�˅��H[J�Y���W�R�_�R=P��L��4HA>c�'?t�φ�Q��ZX��G��f��Oe��hs�1��@�q��Kc���t?M��ڛm���A՜���� R~��Bi��|x)�)�f@��Yv;�֊(]�VPdy��?�У���#�ϝ���u8!���}�\��0����E�Dٱj+H�����p�
�}m���`{}%j&� ���]Ӗ�k4�>f?$�'|��`�7��\Q�� AM�΄�D�H�ru����djs�dՏ�ٯDaQ^��\�E�ڽa�ʜ��@v�EСb��A&�_�!@(��5u�!qp�\��y�fp3iC���^�	�y�f�!�9!���e���	�M����'u�TEOSr,��H!v�6EhB��2� �X��ȉ�Vpg�y����Խa�����&&��yo4��F/�H��H��:��!�K�YW�G)+NP/�N*r䋬�e�����}x�7G�-DH����.��C���^9�({����F��5�kA58m����>�P6�%��h#ľؗ{*޴ekVnlJa�2�ds\+�~��$Tax��K�r��ֹ>�S�@'��-ڽ� �>:�����U�7Al|��ƿf&���$�8*pDr���֜3
����/~�3�Tb��a{��ǆ�� F���:���"�
�*�WVe8�;�suzx�q_��z�}y��l��oj�"�ZPx顂3[ϫ0j��g�;/��f?����soO��]��9�	�4AZG�K�QI�όmE�eA���1�Đ�����%�K�妗�X����[z��s�=��:���.?&j�"��l��C�5�cߛ�� ��r[	�aup�>ݓ>�NǙ�����j�S���'�_+���:�^��_ȷ��c���4��;J�6!ЛڢCx�^H_ʛ��}F����X+#hJ��u� �+/,h�l	�I�	�<��(�|F�̨ �j!��h0�bA1�{��}#�F�]�gg�u]3xJ�1ġ�A�٘4R��ܨN�5�"7�0x��%(׺�r+�\M`"���O�]6c5�B��u�7d	��㺁V.���Ĳi:֋�xlK鹆��6�e*Vu�;�!*�\0t�����]zu0���:��)�tIb�`8�io$9�=��u���קo�xҙB�(o��Ht��:��Q�;Yc٭A��lu]�m��X�<�.U�Z��e���C�+H�V�h_�>T q>iY:�ˈ��3٣���m *�Z2�]Dzʔ�ΧQ��u��@���/��o��������D�O�����;��	� ��j��t��b/����tro�r-sC���eb��=O�J�	D���h��Z��%�LU�?����`��|��,�տ[o��)�Z�2�s58oXi@�uUܹ�7�O�,����e��IXEF�''R�~��T�R�	���yD���L��U�Y�>�][��Q����{�����/b�Ҕ�3tr��o��VȮS,w-��-
�[�Q�cC��l�C��Q�jʳ$Y!&�5wr,�m/���)'�(9dG:m���@_C.epw��Y^�TwX�wń�>�3Eœ��(�����+P���^W@��T̍�y���:��
S���@Я6!L��������WQ��=