XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��, @�����&2�2�����D"0�b�+�<7}ݭ�ԏ�Ź�z�ƋH����-�J�$��Y���L�����x��]#w�G����Q�hyC'<_����8k�E1II�����%r��6��=���3��/Ub ��<	i�ŭh�K���p���P����\|(o@О�n������s���o�xJ�+9�"��fHj�?��e6��%g�T��|߶W�h��g�H/�ݯy�)?�R���.����~4�A�'�o��.�%�;ا���$W����,S�:<�hG�P���Jx/�}>�Fj�A m\ )�v���^�6��A�z���8��s򮜔I�� �p���Ft)J��|Ft	Ym`P:��L�h���˛u���x�IN�gF�Ԁ̧��"x�ϧ�!g��(������� i�C�@o��&�V���-g[�؊m��S��
2�Y%o�g��Ή��?Rh<�����3����C�J�q���5z5�z�P�Xu�+�]T��h��6��<��PJ'�<� s��.ǃ�%���p�U�(^'B��磪{��߽�0\��e��n�Y@n�`��K �߰�J�����+��I*!�)��s��<�Z-��z����)�m�E�3-���@�Y��x���?R[B�;�ؽ����)���v���	���!�K:�й�7��7Q���'S)���Ɯ��BR����YZ�{`�^��e"��*T�U׉z�i��8����i��yk���EeA��<��6=e�XlxVHYEB    4b2a    12e0[}�&O�o�B� T�݇��U1�7�8��J�e��g��Y٪����ox��A�ѫn����f
mW""����E5����G�ڸ]3 �ہߗm�w�2��*�l�Y�[୞�1�5}��X����7�|G4�.�ʎ��I�FCHۉ�F�/(*b6�aB�x�Ol������P'���oJ{�̜/�Z�K���ԉ.[n���8���Ev��Wn-��bP���dC�_~��D����ߑ##�R�XmA%d R���U�r標?39��׶���k��Ǎ!�I�)}~���ЬZ<S��\�'<k���e:P�?0}ɱ��t���md#�=��n��
�/�{;}�D���G�I�w�00��ե=d�R��?k,�9�yr<�$S�)��V-�L,Z�3X3-�'��f�:τ�Q<Ov�_�ӫ#���c�^�ac�^a�����>�hC˼���V�e��ov����U^����Q�zK騔���w�>�m�{�-Z�zd�A��C?9�¥%G肧Z���ls���`�}����0�|ī��xA�^�ho�b�� M�-�P4��<~�1�I�,w,���3tK]
��)��	�À�6�b��'[f�`��Ǣ���zC���޼��%��@��cRq��{n��q|B�T�{n��jq�v?V-,�U�U`!
Z���'ptd���j_��A�OX��{���:y��g`a1Wdch�I'D�p���`�M�N:|���Z0���鑦�f+�@#xCq��L��95�=^R9C�I�M��_d3�����j�>�"e!u(��"w�G_OƋׯ�R8�L�P2C7K��G�G9}�~�z0��9a�0_�wC	���7�^��
+w0�z����}%����9�t�4o��i�cM<^�AY�`�W�$mՍ�(�,����z�$���:�8P�� �����$�1i>�����,�TցO�V�]g������+Nү�����#�D����>lbp�V�|��2�!��IC�8]$i*���U!����$a| �ڞ��W�� ��	Q^_�ێ�$����ޖ��o�{�)D�Z�����q�{���U�*�_���O�m�)��p��F��|����G�P�y\\�0m_���D�"u�\�_�j�Zg]�b��MO+�;����ān&"��
S+h|�|fq�g��5b��0��#���y6˔>s�K��든��C�}��\Β�l:Ce���oU��]t�Jl����?R��|j�$th����GE��7��HT��e��J� �4Ua�-*�ܼ�ծĻ�V@<ey�J���N3K+����New'��'\?�5!�;�#�����,3_���ON��n�0��Y{����Q&�7��a^f&�_��gߕl�|��-�\���1��'s�*��#Šm��'�&s5�c�EA%�Q��ڍ������<��z�Րz�9��|�ĞC�|��
�w���'%������O�dM0~70ȏ�ri�X�ŌѡI����n�@�R�h��m���hb�!�f@�[��n��*'�E��ԒY�iI�׳��Z"`r߈~��<KR�x���1`��Btn����s� I��;�g���o�3�e��%-X��WE�? ����+q�k��^@fY�ri\綛�-}6iQ��"��0� ou�XqI.�4�*�!��];��ୣ,8B7@8�0E0�N=6�-����ͦ�EDƒ�JcM��d#�[��&:5r��~>�>Y�Č���b-�OE��^Sع��O�bm �=�㿳�7��LpK��1zޥY�&l)��uV�&��%pQL$�J�T��)$����s�5N"*(�]b�Z�� ������c���.�Vֱ#Mw�~��b�����T���R�5_��9r��qHk����ƒ*��i#Q��/�177ޤ}Y�jA,���Ĵ:�3�)��m_�u��o|��EAE|&͑__谏'+�̈�g'��g#���%}q_���dy	�l��ϔ��/����m_���:\�)C�N�fݬ(.\&41�Ɖ��P��k����d݀�.[����TX[S�2v/���=8;���/�Y�*�8���A���m���ad��a��Ij��|��!�+�!Sф��2n�>3]�{G�P!���i��4���ąn�����K���/�6�꥙��
�ZX�l�n���	)J?�U�I���)����k�5+���� AX�JP}����%L���
�Lވ���k��N��k-CF��,҄�5l��_M\��<Hp6:����N�]"�`��w���-�'��xt�&(��rȴ��d�]�!�����B��ImA+�S�Oh�ı���W�KDK9xO(�ڦCx�/u� �m{���N]���qչ<�PZ�aٓ_�s�}�H�c�/��3/�SΏ�;k�s�Ԭb��V�v��	�^�/�SG�Y��?;lH�n��B�'�tKn��%d��b4�_=i�Q��d2t����58^I=o�?'y��dA�Đ��ʇ� �������{�\20����!<�[�l}�S��:25��v8�Y!)Tq��C��v�E� "@j��:'Gd��90�Lx�>�� b������A��� D�C���>��<��xM�~F�<���x.?�n��*�{վW�5?Q^,��p%_&�-o*�|���KH�c1�X���/�v��x��V+^C:M�fw�U�0J+z��g-2�S\�A5�*��F���� >\K� >_��"@����r��_�e���-���s���b:��1k�m$U0��?}#ێ˳���|^	MͬA��%Q����'�`��b5:�R�}!�(3�Ć�#�D�ֺ X����$�'�~�23��4n� ���f�\o��`#; �	�4<�N&�I�<�������}�ק�v���.������.*M�E��T��S�&y�p�S��û*[���@w�KIX5ų�*�C��lB�V��3�KB=��&�-����%F鞌�o	8j�|�)�?�A?ja��|�Y~��B�I��5n�� J:�Q��H�2)�[yoj�Xr�*fZ�K�v�b����ֱS>������t�X�b�L�v����.C�G*�z��� OLeXhx��B-�S�����l:}`�hF�\����?��K��)��b� h����RO�=:Km��a���y�WPV*!
�_H�� ��O�r�	��}@0"���0rӹ�GMi2�� ^���>�7�CJi�З����#Pt��N�d W��Sb����;(�z��
�%٥[+$�:�B6~��^hGrΗ�S_h ��Z��<Y4�$Ȓ�x����7a/�Lg���;�ڟD��'��Ifq1!����Z"��6(P��詓���hy�JY��n9U��t�� ጢ�/��邪�0��|U�Nu��m\�c�s\��q�3S�X�_����I�p���>����G�]_9q�E�s�R��id�&�:����|�yӦ$�!����#�1�A5�؇��N؅���}j�#,�L�%UIJq_Y.R �?k� %onK�lE���pP7!���Qu����9�\�I���2	p�zc%�P{�n�;cWݨe�ܦ�38�{�f�>X�v�Zq��?-�S>Xs�h�Ɨ����g-)�KKB��qc�'y��`D��}ͨʍn2X�¦
�{FL��eR*�ӫ���U�:�vk��عS�@e�榝7:�J��a�NO��(��oWO[�L&���&aނ"�x/�2��,�Gs������U���[�?�����8K@��k
F�]�i]�ǴI�Hl�V�$oY��ͱ���N����R{G��Rտ�e��3`�W/D5w^F�t�Qe�O�m �V��e�0����h�>��j��#y�R�p�ȳ�W�$ `�xl�_�ݓ�� ��Kg>��w5�|I�5�<p�nj�FXe����,%��UlX7ƠL�jq6_I�h� <9뽵Q�e�`�^�c
�����;.&�/���h��ΨY��c�|@������a�9����AEȧ�~��6���C\��i�-|=ݴhGvDp�G�
�`��
2p�8�հ�5��n~��O�G�I׆��?�K���9�#*����|��n�@�f��A��O��+	�w����lE��J??�z18I8'�Z����C_1?�_M;␫za����Áu�+'��`��G�з(zqCU'����Ҋ�K/H���z[ѵG/�u�?5�Ɔ�V��Si qh���MDY��"�2����9�pω�W0/؎��9v*_�V�x�4`����f�&�o{�j[������?@*�;<���m����0w��E�����WG�A�٬�D'����+�Յ$�i�!+��Q���eLg�Ǝ��o�p�A�����`�kӁ=W	�1�8o)]���cխ�~���Cc ����+�fe+������Ɲ�tF �"��>����0�Y�@�z�	�o����S_�賁l�B���Z9K��ˇB���ȥQ�I��5Ҹ�+'�ق�f�+��}f��_��������^�i�Eԗ��¿�4��@�7Z�r®��]U��Z��w�$xͧJ?�Z<5/x�MK�����s5e������]B�Zc0�zf>p(�ޗ����������hR\	@X�J1I���Pٍ�4/�m~]\�����=*8!X�K��~��0.#qx�j��ܳ~��E7Ka�Q��� �'�#�ؠV��n;������I^ �1�