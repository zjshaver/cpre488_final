XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����{kҨ?լ�Ő��E�Am�����_k�Bq[ִ��/U�Si����zݽ+�4 PniL'i A�c�`K�r�^QԈ!Pj�O�+:��u�xl6x���	�q���*��gݽ{K���
�#48Qy��~���[;��	�Ge�ݹ�ͳ�(u���bM�>4
@���l�"m�S�d'�;mꡡ`{�����������CQr+CO����Փn�*�x�%��R&�3��Uv�;Z�� +u0�g��J��o�%�˓e}!8��G)v�8F��t(ap^m�(Vm���,����ߡ�a�^�O� 	�Xr�Q����|Q���ΫN�\�N�hė���XMd����^͂Y)�P]ޝK���~ ���^ �F�ފ�p^]d� h��^LbP�=��k��ذ�C�s������������`\�Ԇ<p%��s=3�����V/�UX��e�G'p��P�]R�u�F�ŕw��E�-����c�ﰅ�w�9(�"�7�c�|�²��pI�l V���:b�z�����M��ķ@�B���W�D[���a�ӆ��JaTgG>jz���O|p$)���^�D��x��K-ݥ��H*_�M�U6:�t���q��aO�m�n��c��y�aM�[@AGC=T��5do��ͪ@z|�vQV�j�Ș�V�.X��y�Jv�Tx'j�g��4�|�nS��47���"e9��z�gx�jE�����n�����/��h,�ѫ9�>IȢϿ���������3���Oj������N���R>&��s+�XlxVHYEB    893b    1e30�YBu7��4�@6rjr��Xxbz���U~�b �o�?)�ő���������������`�x
4><S�\����l����ấv*��,]K�f�Z!��I]�o*���.�6�K�����D;ȹ9�k��V�1���f��	{�yuu]d���-�G�>�#�O�&FI��5���f�/��J?�������qX���O���b٭�яX��Q�4+����u���H ���4X�~��
E���M��c��%a��l���X���d�eo7��2qZ\�]�F1W�w��䫺A�Z/j��;���\��&RD%:<'z�,?"Ϲ��_R�eضe�4z+��s�t���m�faN��~����Q3�bǳ�G<��(|�e���S��ի�؜;=SQ�����"E�[>��P�r���F��F�z�|�����d%&���)�g %�;~mi!^Ʒ|q�E<�̔�����:�a	z�9ݘ+�;����#��I��eP�s��6c�ܟM/����>�?{���J�6|����R�sȲ��Yf�W��jQ�]T�z
�I2&r�¨��x
x�@9]:��`P�S������o��h?��M�T��²�J����4걆&�Q\�b������Nf����[gh �T^[��N �@)(�����Bu?�Tzw�{b0:.�m=����5/�K�N	�=�}�#��p�/:�����zV���w|�Hɺ}Z���I-��5)�TY38�j+L�,����7����N4��ML؝j���%����;Ӑ�b��.��&c5���5� �X��`�Ĭ�,�{Ͼ���nf%�E3_�%���c�=��J7L��~ �xv�bh�h�\�Zm�c�����=�].��p݃1�&?�ʐ�����n5�/�
����\q�^L|4�=�����5��ϋ	���Un���B%������Amt�����;@�P@�
)��MTWќ��v+LxmE��6���k&vӪ=/���ԫPhH��]�]���w���&��7I��2*�z��9_�1�\~*�I9�(u�U?l���VRԭR�>�H!��4�J��w�@O�o�L`�5ѿ
�_�������G�G Q+�~J��g;4� ��3��MhU���9�z8g#�0���B?���l�i����6M�����6R��_x�,�`Ul�I�d^`���2���5��w�!D2F�~e��Cy���JsP)�Wk�S�+��`Qo�h��J���wm�M�R�Lgd�ە*>�+��r���w����̲v�ͨ�d������:lc��u��=��H(�Y+�����jǊS�$_��3Ct�g���K+7"�ZE(��7�� ��,�z �d�Ϟ6A9�����X���ü9�#i͍���z���H�
��7�����;k[ö�:Bj�ei�Y>7�`֏���ۛ�Is���>����J�QPE�^�����'�<I�=�prO�����|V��ǅ�d!S���@��Q.��q�X�4�/�F$5�j�|���-���(�W���/g� ��w>���-W�j�ӭ��j;H�xƗ����/��C�zC��{"���B�ʦ�+�;Β�u��ىU��p������R�Kg�E��E:��m��:�+�M?á�:nr39x�`�Ͽ"���`,�<)�*p�d�v��Ɣ����	���M�wj�r�}�Q�CGls]���LWl&w�k�ױ��uW2V^O���R���{����/d�N�l�u�-�|l�swF���-L�]�9���	���b8c���I����*�ے���Ն;M�w# ���c���Miv<�W�7y�>�'�P �=�9�6j����#��j��+F w�%�|�
M��W3Nbcr��,��_?J�~"�I d��#@�@*�O��� ����S0������,�>���g�YXhN�u�[�������yc���j����A���,�e�$%[�h�6��5I܍�����{+�G��[���=�oq,b!��z�^Ճ8��$���}P�^���8��A6M,Uiez�T���W��XP�K�y1�o�q��}��u|�e�8s ���S	��9�˯R����1�xE���ɐ$��Ϭ���$g��̴z5��]h#v��G�JW�%xx���D�������Hnd9Y/���( 4�ued��~L;~��[�t	G��^�3\�|v\�|��&h��TƯc�й�����"Z�M�!s����spׇ��y�������K1�'��=~ ��V0]�+v%�#���q�Q.��<�K٬��k��7Ɩ��sv�5���\��oP+���̾��?>#�L��e�*m0�K.KmY#���K�6y�{�nm���%��N����Q���d.�F�a��u��/�7*0�䝒k���
?���}�2�ČS�f�J=�)�@V�ϳ�A��"4�HW`UҦ�\��������7:%�}~�	"��W�Y5'��t�Yyq���,ŜO�ڏn��� '<�C�{�9�[u٭�|���<]#�$T���d�Z	�0S�F�d�%����c�)HW��ki v��A~�����Il�h@r(KGQ[APݧ��q��.�Ы<�P%���X)(���0�&r �G{����j)_�\Kk�+KC�8���aS&�y��q��g�D�붮��˚�3���-��]��?����!���+��������U&$��~�fT�}uĬ[QQق	1�Mc����{=̕h�M�v}>�'��!���t�rf��̪%�Q�8c��gFV���C���
��l��삪��n�ӧ7%Y@3y�҈M[{QO_$��t�3�e�6*�ѩ�COet�Y�6k��V�b���?x�m��k�L�5H3���W^3�R	���b���*i	1|�K�����jd2�c���Aǃ+��|h%�2ZdH^7d#=V�0	}!n��S��k�.AY�M��ďk	�_�F��` ���dIš5ß��ޓ,5ȸd�$�
֞a2Ln�! ��W}�L�}�`�S4�Γ짎o�� Ħ�W�<
?�鋹H��P�1�ÿy�݊�1S��:��A�$%H��~�ɷv.d��U �-�bVwb�_�}HC��kss��?/���3�:���Ҫ{�8X��1�0�O�!C�-Ң_^�wL$�)ƨ�;�����n�|ӷY��p���̓MUIe�s��u�r8=��kq]⇥�F����v�4����&Nd��B3���P&%�7P��2ٓg=>C=�����n�D#�Lan�w?���88�����C�U6��_2�o�Zj(��{1<w�{پS��3�_�V@�(�T��۾F󃳧6��'���@���\F��'�#K-�,���n�����E����g�D���=��-n�G�@mh�Q0~t�|@� ]�?�*X� >p�)*=��aD�~�QaA�#^����[�3Ƽ^�����q9�G&ZlA�sfC�f�]�l�+g����<�X���M鮞vD��	��>���rҕ4M4|�CϼΠ�ޓ��<mNw��W�4H�p0�3*���x��>���VN���}H�f�k�l�����sB�/��ʹ��]s��q�3kԷ�"l�gu*lI�#�7S�?�̾��Vܫb!��x��%�/��}\K���C=v2t��%[ĸq��`�$��t㪂��ѥѓ����g9�a��	��UM��+E�7o9zʕF�wX�L�I���vƞ8(����u��<%�&�Q�h��v��F^PU���	C���Š+��?|�	}�5,<�;@� �|��_4�X	��0ę#-�eg8Ľ"�$g�{?��}��i֝�,'sn�f�v�Oq쵍"���~:�D/sǁ���8�d���|[K��2��k����o<�z cl���y��4Vkoڈ�4��Y���c���!:�[,����F��G��`HR��Z�"�emY���Q'���2�V�K�y�-��)*}4�g���T~�(xq�4"�0��l�����:3
B�1�m�՗�G�[�����쑅�@ll�'��~�<A5X u�_������DM��O��4#�z�F뱲� 3y&X�X-��6}�f���u�D�'��B9�s���7��)QgY��N�u�/������_��i����:���i�U��V2ͺ2��9���2`�:�w�ꑕ�B��3f��W��q:/��]W�5|;��f�>�7�a�����c�Zn��ki��Ů��6��Q/vx�ɭ�H��qB'^V#jmZZ�3��Q�F�i�Mƨ�.��9��25~�V6c�=��4P����ěFhNm��xW����
����e��Ӵ���:8���p�'�kC�YR=�#Ʋ��h=�RrM�>h��~x<�;���d9���������Q!j�$�ܤI�W�᧳z>iU��j�A:g{�B@5���y�ޠ��i7YQl��"14A�r`��[��DV{���Z\y�c#�yy��5�/�6���Y�G�M
1���]�Z����!1k{�D�"�"�
U.s�>�WbD�f�SA�rN����v���i��B�e������m$rE����\�;a�&��k���c�@a&A ��_A�d�	������?%2&�]]�h��E�Z�۞�b�י��鯋�������n�,Ք=܊���͚G?��[?�Vz��!���Csv�Ie��<�q��/���w_�\N��"]1��R���a���J(&/��Í�)���ۤ�?6�]��D�q'�J���#`�C�� P93��MJ9X�\Õ�J� �Vm�<p(`��N��cfR�q2,,�=�h��&h�Ƽ�>��s2�`�ZzhA�L�9���܀U�A��Z55�З:��KC�UQĢ9��}/`��/����nDW\(?x���哚+n?r?Y�����!"{c4%.h���r��v��<I�X�a�V51���c��Q*:N�-���E��`	O�`�U� ���3�]�|حXU����5꜒tx���!o�^),
�x��Y:��ʯbG�2{i�����+<?�266u�=��K�LlAa��>�g�<%V��z�pnx�\�AAM �A�'2e�ps��y|m��a#"EIH|��b�<��2���U�*f���M@���p\q��S�����O��y�ˏ"$Lm	|o~z��+o��9J6ɦ��ڋ�o1�]�g�vD�!$>���m�)I�d��"$T�}z��}�ʯ��æ�ׅ�S��V4��t�s���|a+����~�=�Ix�{]��dC���wr��+2�^<l�m�d#�΂}��3u�j�p�0�v��X��R�ڊ��'<�D����j9�:~<�4��A;��M3e��{:�.�ޚI?�ʌCU����5�;O!ӏ�G0s>�nχ��	Fr� �~��lX�=��n���*���Y���h�ݘm��~�9~��f��}jN��}y%�O�`�i�Ts�W�L�eA�үB_�R5�h'c�&lt�E�T�M�w�P}JH���o�#J2|-��,;H�H�1����������{�#��]�����V�Z�[	q?��CI��6e*?
�}�"�ܿ�/�^�؇����"�9@�Pn;�&ȕ�q@�'�;i}���Z�����?���* �),�O�P~~�D�~����y����P?���P�{�;������i���dl��eT�A���k���׌��W��]���F���(R���;Z�3�mnB���[>#�Y��0�*[ہ[6����.ӯ|���=Z9���Y���
b�ƏPe߆���{����L�HO3����Ѿ�{o�z�.E����[X�Ťq@��K�?��D3�41,�Z���e�ghɺUկ��S5�����У��쌼������	Aҩ�����(	�������� E��t�u��y��-.�z�Z?����������u��("Q�w�:9�p�|�H����E��zH��f��řN�z�m^��c�!�B�?�G8͐���NO�ɳαZ�!�VBtc�����x�;�iE���,&_S2O81/��:�����a��b*����RQr�8�:�������/x�	��)�/f䈏��v~a�ç���Ρu�~��b�Sx���%�}8�!FT�5΅�')�y ���,� ��pK�_l��A���_��i��5c~o�R�P�;+�4ة�V�9<�$�C�w�}k[���\��}h�ƍW���a��O�<_�E�{�X_��n��8}�.ɣ�)��*��XRĆ紒�.$8O^�5��)Ls��$�謧�f
6���ar��(<��FC9�����V�
,�)|��:�����o�����|O����f�B��p���+;��)��;q����w�>c� �͓a��cW����@k��r��bqr�B�ЏܶY&�O��r7$�QX佶��v��腖<\�-G7��f��B͡�}��=�:x��+9���.�_7�;�V�6�C���2����J� ~obf��P����P�O{��@u��4r3�⢑G����r�>��Ο�Y��Z%f����ͷ\�Qݚd~�����S�,�Dn0���i����8C\4�"���>*V���f�	k�1�]��,���bŋ����s�1�9.K}�@�.�٬���S��+
Т�V1���i���Z�863����)���Zw�u��B0�7�q5����Cr�:���$��<i�P��[�wϾ.�<�a� ����̶z;�VTq��J'�C��T};yy��$��>�p���H�E�ܾW�i�뷤 ��/Uʴ����8#�\�����{-�A��@u]�T��N?G��D�:�;z��S�c�ep���J�0���(�x��R�l^�pϮB�r�7������Kdq`/�F��J\5�;3��[Z@��\0L����Q� �!�%�J�c�G��{���X���eTU&x�@�0�16�L��v懜?q�t�'�P-�l!��Q���=�H?3���
½�q�?�l�&794k�'�]�н���F�3XQX����SyG�]��M.�������Cq���?d����n��$	�E?V�	1l���KS�;�T�@y<h5p/���8W����g���ʍ:���roT�bQN�U�Miuu�ާ���$�I]|��H�o�,Z�V<_7-�R!ki�n�w��1���eY_�@٠>�ƅFIo�/�6�?.J�;Y�
fs�����\��*[s�q�����n�o�P:w#��V����-��~��O=آ����[>�̦��g�n�j^�2��� Z[\�w��]��M�>�o)Z��r��6^������CD�.O@Uͅ"��X���w)ܮ;9Ә����Rs��5��uyE�U�W�
^�D!�������M�?B,�n5�C�N�1��&B���s��(+u��A[��w,���3l2�]kݭ�'+f�E�~��įL]p�I��Qv� �z���kS�n�)��"�۴חʿ)H|�ZSY�i[�#��F��pq�cI�uu��(ص����~+jw��_N��nk�R��nޞe	��R)fJ$�4s���,Yp�'�EE�*�"�h��ѱsb����bi�����
!�e�fJ:��'�Hۖ���k {�&����U�j��)�