XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��MC?rq�m>��o� 4�_2���;�/�׾��qxE�&����@ʶq��|�_so�w	F��K��=�;�d��:�/��Iu*�0�O�a�,��Z����=Q�b7���K�n���;��v�n�{�!¢'��4wF�g�aw8G׍5�M��S=]y�Bd�$�;�UD�!g�,wqt�
v�O��ǖҙȒe�S=�����^���dy�C��D���u���EP���4��|D:�*_<�'!/o+�*N�+�z��X�Y��b�F5N��Ĥhr�hQs
�A�C"I�y>Mv��#���&jo�9)<-�8@���F�PE�`mn�~�6V�t7�_Z�e���'��Lh��!���*��EU�ܱ�ŝN 7R�v_��I���G#[��U�m�$�G�q�Iz�S��xOyF�.h����:���5�Ѝ���) ޖ�P�3�2�l'}�$�Ԩ�����|E�wP���(�|9Ȣ���:��*i���������v"�D��!������<A��%ɖu"�~	0�d-���w�$�.�6P^pDY��s�j��jP��$]��ұ'�4!���A�J'��l�ϿU�x�����k�>�=��0��|��a>�� {���r��k�)�I�|�_s&�M�A^3,;�Xs�殸 ������^o;v��Q�����Q�v[qW��X�aD��?�͵�٥C�6���-Ҹk̃5��ew��Qo��e��N��I�$K���b��0�mZ[�Љ�����sj��XlxVHYEB    2326     980�sW��녅,!�!-�)P�6�w�4�lH�/�a$]�0�S&���ĳ-�'���7_��$r��wa���u@��I�����o���.�w����l1�'0�Mg�\S:k��ǚ�m�$C��r�\a��*����},����m��]�\�|M�˗PP�JA��U+����#j,�gU��e��������Ayw��|����k��O�N�K�lj#�̽8̋.$�j�*�����}�w��D����g`H��!Z}��j���4�(��c�]�9Z�B~�V�O���W��k��<����}Zg4܇ƛf�0���2>͢�k��C�Q�A�,'�-�o�t�8o�P��[N�e��{�:T*���c`�L� ��:VPR��3��-�]��ZT���F PA�:Hv:Kk@��ק5�yO~R�G�1>I��J�x/D	K>Fd����J&G��v6�� =����l'k��W�����]�	����I�����tp�J�]{绁q��Y�:��о\厡ͮ�S}y+%�������d�Ѷ���,��7I�6a����
e�~_��rͬw�H���6�0�ʳ�~�d�M=��P
�l������;8����<�]�Z2a�굫���i�t���r�a��뛔ٹG��a���!��o�����#�����pFz�YxЉ���s&�@,�%�D\���5��sUB�8��s�2��!���6�rk��×0>��������M�xBK�F�, ����j����ÜжrҝLx��ݟJ��@�S��Q�i��c���u�8L*\�O�o#��.�+6��p�>�"9Z�l/c�]�;P!s�i�����ǹl���d�N��7���NE�HJ��k$�_�ckxkiF� ��-V��݀b/(�
��Oy׶dmֽl�`�#Y��fH:�ʟ@���<��4��05k�L�KM$c�Q�:���w�ƍ�STC�}��L��_�5����R��yyQ��2��6���`Z��\><ڦ�Er،p�&)���m��R@�Ԙ��s�)�}r+�#��=yD];�Q���Y|>��J��6yd���>���n~�n���G9<D��X n��T��M���J`�1����s�O������J�h�:�#@R�ߥCK%f�>��=�'̴�Q����htRf%/>�.'.�W�(q�$��g .��pe!��D�윎�֝l4�KZoĹS��0�ɇᬞ��_x�Y���y
-TϚ	�T)�|z� ,��(�:�I%*4��kGAB|#ִZ�۲5��j�f�#�QT�Z�<<z���K��c0VȳcW�K�>|�h@ ⓛ�j�,����]	���w��Iﶆ�*�h��3 ���ft���\��|p��A)����.�z��Ѝ������
�L��	 �,��@K�_�x�r�[���?�,?��=��\FgO5y���Hm�}�qp�ܣs�j�ݞ�@�`�IA�;^�X&���ЧR�B��E`R��Hd
�4�(Y;�#�7��N�ҸAXSTU�I�d�p�'(vW�4��V� ���f��y�����}�C�}������P꫷kI1�����B�>�(��=+�e;��RA|X�����H�͖ƖN���rd��@��q�0c�_1�_G0Ծ�;g%��0�D=��T��r��b�>�<<T��)������I,A��Zr��0-7����>�[���7��T�M�>�r�2�Z�<F�F���8����S$52/���\���9|g�����-��2ՔX�6��+�����/
���.��6vCT���qq��u�,�I�=Ū"����� �/��g�gZ�"���p�h؎Sbh��h�G+�%�X�qgb&��H�&j�.�*��K��g�M��5���" �]��'�&�������a��X��9��樝M�����>�������Q�!��n���~��'��7��va|[E�Pu�� icI��T���S4�}��RV
/�
��O�ߑ@�� �?|#�6S�Z�Ԣ�\�s��Z�jx<�M��}ն���%ɳQ*/�t%$�l)����_V�~OF� fP�ɣ�+�X�
�I����#�}��`���b�ٱ!P�̭eB&�dϑ��M
�ʖCAA� �>���D!��\؛�6WCRH5��+����z�I�Z�1���P�®pB-�����g���k�8<�졇i㧌]f�e�w�Z�H�
����. R�6��u�y�-��X���j[���^;�;�zq��Zٳ U�*`�m|,�#�D�\+N�]�e��/舱�|�ǫ�Iŉ�_���Gqo� :���\����1d#X����j��Sy�W?�c�-���c����[n���Wg��br)= -�\����<z��h���̶�8>UO{��