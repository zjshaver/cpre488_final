XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��]�B+3���sE0���'б6hO���/�x߫�mZ�z�'�vz
|���S���o7��+�us:@`\>���(<y���&5D���������`a���&�y�K�5P&���i�E#+8C��k�����x�>��{���+�ݴQ��
T���Cɑ�+au�3\ѷOu�����eV��g���3�.��Z����8�8�/���No1u����ᳯ^�&������P�f�byvX�<G�A�j�[t�]��0r�4;�=9�׸%�
���@������[��{�?�ߝ�+V6@r5W�x�Qa/�? 
��_�
j}����c�+�yLE�����fp�
i*or��><���$�T��>��/�V�S'��㥑��n4�m��<�Sn��@�=�
�p�A����x��B�	�ׯ��0��������������\ר�%R�l�*�ܖ����
0.�@�G�z�>HGπNHS~i@n���YV�'~\;�r����ϖV"}?�!pw�.�@8ūpG���t/@=j�����X��Ƞ���,-���	�
N[��D���a�V���r�bu,3�ѡ���T H����(�GI������ǔ5v���Z��/.��D��݊w�Z]e�k�gx�
$�ڊ4�Ń�_F�+ۿ |�0R���@���\/*�6?��?�VgV�? 	���-�R���u�y�&���?�&���q�5�t�g�ݙ@�XlxVHYEB    241a     ad0�&�~�v���ѷ׵jtn�'(�aJ�_G3����a@�tЎx� �cp�����+7Լ�|�����Ņ��bN��ķ!oI��Z6x}�<��C_�8̟���ȔsT����g�_x�^�Nc�sl++9�Fs�����On%M�m<��׆�J�*VP'�	�����c���x�Ƽ^��译DMr�5{��K�ck�/���4i����|���wѨe
�x��5��:%>;>��N"�_���PQx*SmLP�2���Ʀ��Ub�d��^-Y�㑹?O@�;ǁ�5tbsqq?r,r9�;�,y�E'��a��S�>C^�,�Y��Q2P�#�����-ԅ�mDsu�),|�t�9�K����ԸV��pN�܀�nfgM�$ڟ��I�jc�<��/`�1[�GN�Vq������>yk�ēw�%~V��Z汄��P¶�1����"�L�B��?�5Ԁ,��Tْ����x�J8yl�<���i���#nu�x*2I0vOM�����z��ą`���U�i���Mq��T�̃A�ʐ襦v�@�0�^c�ܙp�����6���?�fU�d�����V�yG���QI���K�	c%����\6:y>�q	���>@_6��ă"pºo��TL~������y��p�r��C���9����г1����/��Lx��5�ӗ�nk�UW�Fe
To{f֡�y���;x�S��z�ΟY��o`Zo��(����B�|�]��x���_�v�i@�6�]�aɖY�EM-�\=��&�����x�2���ˡ��$�$�'��gm6�qc�Xz�O7���"�]x�O�_���ħ�V���QM-z�0��=?�O����=��f�l8X�:���O�_�N)�Ex=��?2w5E}uX/�V��P��? �{ߖ�a��;�.�D��{���)��=��<P��zP�6֙1�s�`ٝ"T�Z��p�k��.�أ,}'[�K�~U-*~L=��g 7b�m��$��ʲ`����0P��������n�7�����#@��)�aq�,�4ih��L��1y���B�,�6�âI{��E���9���V���7AW�3����(P��'۰9���	��i�c_����qϖ�I�)c���M�y�@l�毐[���4)�ޟݣ�a գ��č	�>Z�]��n7��kNi�zX�#�Fsb_x=�vo6$ݤ���U��.�^�����t�W���>ӱO� �>ϙLE&����J��`�"�I��cu�p�����ˡ�:�4�.?��o:Da<�J��Dv�O�y���+�����^i�~Z����/r^����[k��%��r����S�$��G:�R���ID��pm���u� �ĩ#c��d3��_���κ1�U��҈OP�2�LE1k>�k�/��O�k��~�nQh����r��A�z�y 	�c��Ǹ��∴���31ߺOa ���&����s��wkh1Wy�7Uv�9��B�o i� �$f]?ܬ�P��3�=��A�/9%g��ȱ��B���a�|n?�N#pcSd^6q�?�d4\;ZA�;I�O^@�|j�^�l�Y�cJ7	�%��v���!X� ���&VL��5|]�Ry@�L3����48���,��a(��ɷ=񍕖Ȳ�a$.�1|�+9zlh�+S���W��*�߿�����B5������Gp�ˀ}Wq��D曌�[���?v�A�%��P��Ģ���A/I��n�=��Y��>h.cBF��:l(�2�L]����ܣ�ƃB��P��+�k2��*��]���� �v��C��Ŝ���� �%��~�5kY�Rj�=����	�9���\�?R�0��Y�d�~'�!"RJ����F�$D�з�щ�K����7��3��y}ǿ45�j�W�:�(�@L��liW��`?�V�<5�7�� �5_��ێN�2�A,�0>�YFl�w����ߪy���e��D�eO�ueW���K7DM5��3</'�;� Z1�����p��i���*Y�����_5�����Y4Z�^.��L�5�3�;K�@u��r|-���Dvf�k�/��F�+�Xm86i��"���/ʀ��Y��b�1�]HQɡ����9��GU�J(�lS�Q,q�lWTn���M�g~.�=��y���%�ֿSY�	z��?��إ�N��Rh_�&O��䤧��A�r�?AHp"K��Y=k�£��{��-��L���S���F1l�x���~��@�(��wմ��B��j���X���ҝ�䨞8�8t"V�y�D�������sZs��y��/���w�z���Q��꧿����w�+
 ��e������b��U*�}��Yh^wv�N�F�8��X�Bޢ_��%u����9x��C��2�p-��f?����'+^�'�%��� �X0�Y�\���5Ϊ�:�6+~�����i��f�"�8�s1���4Ih�C��^l8�v�0$n�����	�Lj�t/���k�AWz�����1_���̅n����b�prĻ�o��̄[{����@�;�՜U�,�n.
Y�7�`5��;�ϡL�4��L�W?������SH�V%�z�-&��w�_;�2�~�w��&QN��E����_���ŷX��l���k��b�I-4�N�����u��+R����=>�-$*�0�/��,4�A�ÏjJ⾼���b����$Z����