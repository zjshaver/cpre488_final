XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���G؅�s��f��3��Y-�Y�wk1���
��-���)�Z�fƥ��W��A�R�kˈ����&�RkХ�ir�J�X���a���N��VeGНM�b���Z߉]�qK�""5N~daQL")���o�����&D�T\�����o6�H�>NeO�}�W���c�����s��OR���@/���l�,��k�Wa78�����Ä�s�DpP���s�����U�HoWV�b����C&�~�|k��xE:�2�A�2�\�Gl�rN�3��`t�w�c�E~9�#2���w��\�~L��z��lЊˍ��H��]����q�ń����M6���,�uԯX4��RJ�*H�ݷ��
/c6/�w~���*����:`�$���
�a��µ��M˴/�H�~>�d�����^�΀x';{�Qc�bFw��H�H�-`�QL���M���Œ<�0પ�����A�����
ɝqn Y�^�є����B��5�-�:���6����8F]�&M�*wf:G3�]�F���1�e��؍�筇l&�A���"ޓ����d���N�2�U�z礥�ƈ��VJ�n�t�f�m��Ӟ�h�>}��Z@�!g��L@v�M�!��|���:��L��P!�,,m�_o� 49CF�8O*�sF��_,"{� ��x�� X�����C~臡���N��_#��\�28wl:ߦg�`�KO4v�d��i*��b�W���s��qB��+z�I�XlxVHYEB    af58    1ac0�?"��.���!GZd�F��7l�m�7g�D7���+<����6��[�t?��H���W2asV���M�`�x�V�ː%+z�H��N�|���?��'�_��s�z�{���jB�d�Օ5�8��c#ǵ����Z賕�H ��~���r%v3�j�Q�
�B���&��Z�.���y	ǅp���tK<ٕW����P���wY ��f���C5ńH:I�h"�� �J��{E��x�+�6)�!sYNd�ĸm��� .��2�|�(f��w��q�eJ���DI����#Bt��-��P�<7#F��d���)+Um�~>�U�\��Υn�G��>~��9��B��[G�))Zr)�7���ŚN������1r�R !��NU�s`6��7���FE������ܲ���6Z,%3qV\38� ��M�O3�$+dʦ9� ��^q����x ��d���Z� W��A3��sd����?n���J��J��]�s�Eʃ���㚹�.�t��.#U�C$�4��h�>e]��^d��k�Nb����b&9-��A�K��+����J}c�ݒ��mi��<���Uo¤���H��������70sZC�=�/�_D��@�K����G�lV���YIF t|F4��<��m�m�-3�"����r���9�d������YE���d726=���B�8��5J@g()�HU*m�/ԋ�\aP;�;�h���|8��}M�R�S�0����������;+�%�	ׯ�C�tR D��1Ӑ��~������4�&��,ڃ�&AY�-��6�b�pJ���:zD��<Ͳ噇��Hh�5F��0=Y!ri�v�B5j�mŔ\�>�C��Y��J�~�ú$���7�3�U^U���Σ/�96��7�p~���^,&��m<W������%�(�ת�(�J���mƨjՓb�g���.��1��]);�*A=���(h��Upu��IK~䇵�'��)��}��Ѻ�����#U��,��%�w�Sn��;S\lb��P?Q�..#N�c�JS� �)p�8�F�:G��6
�"AT�W
Eb����fh$<n�ⱱ�U���Za�߆��K���?�1<�o��06BϢ����,�W��\���!g�+;��kdN��� �>nG8�����,��6Z]�]�v\��_��,��Hg'V4�me`VS�%:s��t��6 �X���M���#>.eP�7�����{�8�ǭ�1����X�� ә��[�J�;���?Lg#�T�ʛ'Hj?V=��4n��kv�{��+��R��O�g��8z����"�4��T��8�#	�Y�p�	����sq��Q���V�V�̹�5����(��W���&�3�:ĥ�/5ap���(��u�G*�?T��1��_G���+t+����S+�p�IG[SxA����:��Mƻ�:�д���4�S����f#����!W�����*�];v#�W�;�3nk,�!͌�*ې�I�m$��7#2�*��������������Z;*>�}��Ry��ĉ;� ����q�`!����q^�
`��"���#�X���
�q~�|��6�T�dC��5;�%P�|�h�z׹Yﻹiu��~�v;!�fXuIVӓy��Eyn��O�����|�[8�EV뱢6-k%���0��7_3��Md��B���
�NBb��KK�AZI|�%���G:�Ů�����i��8��'w�eE�뚍][��p�5��N�A��h��DM��o�(�=�z����R9��;q�u)��l5�5����n�>{wO��L�����m&T�G��I�7bH�0[fh�1�R��r!��@&s�/��ݤ�����ӌ��yˍ��N��ܬ�	�p��?u@	^�:�O㢧�~KkTy�Ѓ/칵G������W^�	��`�{��q-��(UbNi`ms��ͣ�c��9���#\���N�ΗN��j/⥻5p ��!��^���?{d�T��?�!�r8X��{i��i��� �w�
�H�8�ĺx�ϓ�s��D����{'��d-�S�U|]r'_����S�揎�0��Y D�����ǵ���`C' %&��-q��6�7k��ƳA�����7(&<��CJ�Up���v�Z���4��<���E���O�Y��]�+��jZ��T�}��콱���Ĳ8��@�ae�NM�½o���|]!���OvL�8+
?��7�[��uſ�F�r��z�[1[����XjD_gA���Z��E�� k��� *�nh��Xb(>a*�	~������y1_֊y�A���	���j1.�;D�K��X+r�������ߴ����A��=�Y�	#��A�ӛ�d��rTW#�e˩�W�@:~���)r���b2b��K���m-��z�Pu�1�p����Nz����G`m�"j���H"�%��.qq��;;�Oo�o�X��Ɨb ࡟�\V�����h�r�z�_��ı���x��nl�ʹ�3�`oL�m%���n�g1�� ���W�\r��3)����@��0���=����zZ���.`��K_���3?�z�${83݆U�N�@�~i�r�?�:`�3/`R/��c!?��6���M����ɮy���Ipٷ)
����o%��N�ch�ҢN ���[���v�rJ�ཪ�i��$��5�������M��FF��ܛ،L��}��9�R^W��zx?��32��E*ѵ=����hk���30�}���O:�P��D�Ύ��(��A��Z/����;�ryR��hV�mW) 9���S/�9#�S2�Ժ&S�Wd��*]��I��aX�W3��|�Ο�>��C�:r�̧����Va)s���@0aSB-_2��/>�H�eH�L�S�E�?�_��f�b���WjUv�J(ɱ�&��M�]&M��bT,+m��S�_\���a�B�l�0�h�v�����̬"H��^v�{,.fD��H|%ݝdm{Ҡ,�v
`	���;�YJ����E�8a�`�IJ�3e�K���S���R9�3҆~m��r�	��|@�������i2 �Cr�'%���y�������5	��z�c;���ʿ�*<�uPdP�.�5���"+��A�����}�$���%ߔ�:>��B�<��� �^4���Zؑ�ۑvN�V���4�Ez7��]Ցc>��x���D��tDG������V��~PB��m����S���!s�O������l�r��N�H�0�\\�9g�\*�Ë�6d�˩�W�ZwO,=5_��i.1,6�9nԼL�q �y��m���X0PO�f�z�GF�Ƥ"��5���)��c�z�՘6t��8�)��c6��)�8 �;��Y������8FL`�X�bZ:yП�)_��%i���~�7́�A:Ek){����!��.�G�kUf�(�戙T���Sj�L�M�b��Ϛ����vG��G�m�i���x�uBi��u#��}Ar�#O�=��b4��H*�1Gѫ�gZ��Q4�:�F��,�q)������e/��Jf�M^���"�B��䌂�P)��}��067��=�$eh=OՐBQ^��d�����7[j��8�s�ǈ:[�>$y��\�O�ڂ��S�v�������֫��m��w��P��8;� �]���$f�b����}!���q|��K��s%��8dz:!Q˥1�#���//019��A��T�ٌg7��:��E���y���W�3�����3hI!~�~*��I���z̸-6�&1O����W��8+x'��T/b�u_1W/	�A�ʊd��({�SՐ,2܃"6����ʙ��K̢�`��>T�A�Ժ�� M����c7�o�2�cל����%��G��#P��6��4#G�S�+TQl���/�rL8�m��;�f�Lq�n�i�28V�P3�ֆߤ[��P9>%���m��M����Z�Џ_^tu��q���w�����?�WŬ��4�U�����0j�#��q��h�:֘�ΰ�k�3��}}�R�5������F�"|��u��E
�N�l;=�|i�&ѡ�к��X��2�MP��Gc|߇l�s*�4gsɁ��/���i��A��%�}`��)0��+��feN�Z%Y2�e��?��/���G^˴X�g�+@)����tB�NԆ���*�QX��[k�B~�~IT�=�qV�K��-�� �NƵ��"�{�[�E
 �ڐ^�jZ�ތY�!�hѝ��hv�r7�����mH]δ����bb��Y�Ȕ񦪍�Y�n\s���o��g+�$L�?w�)Y��(�B�8���g~������k�l�h�l��pP�<[�ޡ��0��F����BU}����d�`�$3��Av1U�qU��)s���G"� Xuf��ӵ\�
r� �iR��Qg9|+�|��
�ך�K�t��Xr�6�x�,��r�
�bh�p�չ� 혣1	S��m;�z!bd99)s�d
�Ķs�Y��ESh)��z�f��9�����?�4�)���f�@~��.XLsr>P;׆���<#�Z��,45;u�P��-�����Vс����� r�����Ť�z2�x9�����9B[/���@�I�`E��IPc�n*B }�	��6��?�f)�A�_t��+$�􌑸�fE��E��#��Z���U�ܗٺ���X��x`�Ed�(�O�i�q�H^�p�va����i�;�p�bX��<2�5�b�}3�g�t�p,K��2ƥ�u�PR��a7P� �����S؅�唟
)��U��]%$؊H:�6~��ȷ�%��r���ꌣ��Xy�)N�QPN&�}��3��J��
2�^��rz<]�̼����W�a�wy���\1ҩ�U����r�^��Iie����5	�!4/YL��;1QM}��O]�s�R��eF�˶6�Z�)�W�KΓ��X~[.��6އچ	�\
�}N�GP�Ɔ<��/����y{������ؐ H!yVf�-#vZ��la�����!���3an����G��q�ݙ�r�d�'wH>Y);�K:2*�]�a�����
L=jم�ΜW���wQ���.Z�L�Bi��^�=~`���<>��2�{k��G/�k���MԦ�:u�X���;˵amf�]��.qBF���[���%���In���F��52��E�	��<MY�4Ǝ�����4�l�P�,g7G{W��S,���E~�;�"q>k|�"wބ�f�\�'��^�������h�0�$,������Iv�DG��.��ӑ���U���������ͩ�舒�.���t���n`��H}�(J�������j:�{��]J�dN�~5�����O@;ܼ}���7���HY�>��"���@���G���ڔ�[rOH����#�����Y��A�90w�<Z�k�qmw"�V�NXFR��A�kr����4��_�|9��n�6�Y��NK���9�k�������&9�l��z��$N�'�ʊo>�Ɓ�{�!�\��xd=��`��E�-:��"tp�;UA�U�k�?䰀�(��2"���*O5&�=#�T` S��q*e�;;����pMڍ�]�u%�2���ع���x��.M��Z|n�u':R���r��1]z�f�c��Q��wp�-�
����^����� 1��o!��d �~�J�y��˜��B�M����9�E��b�e��F H��k���C�!'c��3Kz�jBm�V�@-��A��	$��X�Rj��W�(�#�ߴC�]�oM�sbG?���ljp�aP�&��'��c����Y�/%�M@�b}����D�>�}���Oڂf�r�P�sc	�[�R��+�p�b��YnJ>2{L�SR���������й��.��7�Օn=��c�5(K�B�����i��`M�6�Ík�ÕR���Z��Y�1���N` 5�2B��f���\�w6�������3_���H�]}	��	�|N����ܭ8�AEe)ҋ����*:�xlf<̇����E�z��.����� ���`�^�M�?��#c�&�\rᴵt"�po��H�1����M]��A�Cb	�>���&�������ٟ���+�j���Sx�*����ģ�������0���9��󧣪��0�n�~��S|&�U��S��Cߍz�>JB���<�Vρ7������v~c�#�޻Z�y��=Wz)*bwB�����Km�����:w�	��l>VF^�(U���&[�X�g)�k�t	{r���(�,��h�;}�n"�cZNM_����P����"�P�
#듾F��^�M��QShMz>){��I��7�A��m؅.ϲ]�؎����?���z��@�r�L��k��mm
�ft*�1C����jڸԴ�[�ʟ��k�64�D4��n�$�ň�y�u�W��\���%�u�:ͤՙ������@ V�ٟZ�&��"����{~\~{�2��� ��;x�~�I�������(�MX ����>i��Z7�93!f�A<3�.>����/l5�kg�s�h��qM�%j�~��4���9~�3�=���)6�=۞�2��r�E`�w����꯾�+~��I%�@/@xaziΏ���{�cE�a�p�뤩�V�h��Vv�Y6蘼f�4V��	N�ɱD�Ca����5VQ��ѦC��{���yT-3�Ჩ��F{#`T��