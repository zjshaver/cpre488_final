XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���7'�\N	Nk����@��v��A�@.���	��xj,p|�H�ꅔZ�����t�2�;Xj��XԞ�]뜦� ?i��|�|��3�6�=��[|������`�Ԕ�G���&�+"�`�`�����<��}�x����$b���EXJa$�;f��I��褮���u0}txk����|�,�W�+P�� ��W�ݽ���1K���V�z��{G2�w��*{
������>�S�2�}��/�&³k�%�$r�Ӵw���:��Y�q���=%^ʏ9�hѷx��u��fn�� �Y�-W0+'5;���W�Q�sj<g�֥#�2u��yzKV�4cp��m+/�謕%8�����,�����}TV�cr��8�{ _�W�L��	{�5�:�q�w|�
�}�'Z	d��+�h�C�_Cl��<��;���՟g�0�vl�\�k�5��}�
��ҁ�p]i��O-F�Q�w�`�SՊ�\E ���1Vu~���2i\�\��c��B�w,_Ef�l��l�ARO϶�fr�(�� r��.�Jʂ�}0�d��	�Z4Ԃa���^����7�j�����μG��{n�+�4�x{#KN��;�Ȇ�?�c#��DTc6�ul�#��[9JfY�)�@�U=�	O�f]��d*E��w�����H�E��͌}.oܗߍ>��!�)�������%#�!/����Cahz�]�pO
{�ť�v�>���,�m�k���L�yqXlxVHYEB    2b75     cd0����>�xo-껻��a�
Q�;�Â����xo��h�w彛$�)&�=S���J��`s��:�b�I�n+X��E�	^�O���}F�m���`:`�4�Ǳ�(;Ү#.r�T��ܙ.[�h�X���a��bO�� ��-��m%<m_8���ݢ����`c*gI�V�U;+����*�i��U�=�FO����!4c��q��C΁������y�=E���0֙�.�������M	���>�X�+l���k��Kv�z�>v� Qot��i"����bL�n ,j����ݍ�/�+V�/w�Z��A`��}�� 6�Ҡ��r!�|��G�D^�����b�褆�b��w�|� �Wɺ���U���v?w!!��%,>��,-���U"&�����ÿФ(�XX+�������P����J�"�,�}e����d/�P.��d���!;��FȰ�܈v�]��k�e^RO�2J����m������'4��ò�3Q:�3;��Hp)M��G�*��:y(96��v�6L!}ʿ&>��-�)g �0+��Ŝ"$P�X88�Y߾G��7�D��$ј�J�݈}ilW� p%8���ot�
�Yz9t���'b�|���>ؐ�88�H�HQs+�����CG�{�(
��o�%�!$R�T���\�5m�����~���/$Q28QШ��|\�ݠh.n�/�E])��yth�t��f�wXL�K�v	��bUaC,_p���D�Ҟ��	��G^ #	�m"W���?5��5aEY`C�evTnr�M�s
O�����;�Ի �&����WM�R!���Mm�E�X�*�ˎ}uMH|��G��+�����e�֙�"!uq�8Q/s�<�b����׫�~�鳅1�^�D��'�)�쵟��)���
P4�J���Jh�WT��6� �O�@S��c���$xUgi�qCX�1~N���50��**
ܛ'��??i��0R��N�	�Q��]�(º��]�z�����6� �J�����A�1O�i�@��FC�1��Lqe�\�V�zH!{Dܒ4T9�V�����˴1u�JE6�c�o⢹�Ĭ�7�O��}�F�
~9 �"�����4G;;}Ѡ?���sY�eƾL��5-��ݚ���X��D�7��m,&6��-#�?[<x����6m+I����FIHz�}Ԋyt�;!阓�����"�^�/����&/\�'�,�2�n�ٵv��C��%꽞�*�B��ݞ"r�Lg5H�����k��d�$��_�Z��c�ډ��d���f֐�զ��@{�K��nU��}Z*�w�?�ݍ.@E��Ҩ�7�&��`B%,��~�E�J3E�Fi{6!i"QbQ�Fx<V�˰u��[�.�G9�~셌��W���GuI��n�c��^�	!R��<nr۴�,k��R�X�`���x5�xp)�������ntܓ<�U_x.k1�ݴP��3�xV�濎`��{*��O@��&��E�*9Ç������Sk%�X��[����TcF��6���Lw
9�2�8~�a,gpr`6�E5����
�����2�Q��	�c<���U�#��v�C0s`m6ػ���6g^�R�������Ƌ�\�%'���\.�-1��pE,DU�0���|fWI�g���<}�1<�5�c�g�Lpxj��:��T>����[�y�%�^��T\t�{�1M������C0�#��f�]�m���z�Spe��<��27&:��Z�v�� �M!/�1y�Q9��c9	b<N�;�ne�K��&�C)�9l�|}�&r�.$�z13O�T��:-[�͙��u(��^��|m�� |���nI�e<���V�Ԭ��?,l�f*_�c=�"R�r_�i_]�I��mu���ߟ	��T��P��m��S(�����E`ϩ�6٣��i��9ۿ�$�����@s�1�8ky��޶��)���%���y�KwG�q-��o8��y�L����Ҙs�#������<O�/����X>����T�� �H��ګ�*TN�/�&��|;s���!�E�id�T�[��I��ζA"�O�{\g�v%8.'!�����q� ���O!�=�G����ZN@x��@�6*O��3Y�+=!�"�������GC�B��G
뷱����.�<�
o���h-�d����s�J������6�;�i=o�;���Q �� �iN�=3E
7�2�\~(���%a�I�D��F��qL �P�o��1�<"\j�����}�0�IB?���2�	�ߝ�\�(�3|��K�#?y��##��߫�e�{;��'�sjɬ��2˦0���]�Zq$s��R�{[�݊:�A�t����?֋�J#�<8���6�����j|X�����;S='kM�h���a��hw�����6���;[���`���������x�!��+cXp�d���Иo�[JĮ�0J�z �/a����YO�����'�7�՝U�7 ����(��}w��Et�2D8#w��W#C�z�P뭄�4YM|l���0��E�e��
��5i�+��+��EY~�H��T;�z�YksU�A|��$\mI�_���el��+��WX[&:ύ��ɯU��c��C�n�xI�2a�P��S���J���\��׿ N��M�.��dݼ��'	�w�W˯���-ͽ��h҇n��	f]�X
�ef����Jq9��.� &�-�1���.�"b�����:h1�w�i(����>:��1�m�9Hʾ��`���h���g~��&`���@د��g��Y�a���r���F\�6���0Um-���Kh�P�J*G��MPd+�!lZdm����Pqn^�]�e��(�����J��>����ԄPz�5~K�FХ��3R�'�+%aH{N�]4P)*MX*�&Uq���i�� ��I�p@ ��^, 	h���Sc�9���(Da�3<�3%x?�ee&i�
%�ֱс0���Gf�#3���x�6�
�O
cs����3v�]#��z�f3���sgG�؟��-�����\�2�˕�Q�e���j�����[�ˎ�J�̾��$_�k��rԱ��/�t�yF �z�m��-���B��}��F��ܘB@���}���#��9��3����5���WfT'	gl��=���&h�Ж�5J�Č�H��O!���1A>Xp�D���g� �Ý��--��h��k��,��Ux�