XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���mme���8�{k<>{Q�!�{�t3�;�`�[x"� W�ã��*ƴ$��z��J��Me[ԅH�횝��&RG@k�F��]�`�NF4�4�@�p��[���0��:��P���ds�ŕ�k)J��6�dy g����/y����"�G ��_���ͷ�ڐ�^���<W�=W�+�|lVq|�f�,��Mv!av(��K~�mV��ڰ�O�̈�n��_6xn0���*��MD,ȪL�֭�r�^��>��nL& Վm��/Б���z�u�E��?L,R�uǊ�m��Ɍ��#���/%��\=gI���;����%����e42Q,ؽ���B���}c7�at�:p"�Q�NHS��J�k�(��Q�O�|���Ld����V}�h�\45F�>���3_N儺G���Xa�Z]#�f_s�j:�����z���wߍ��v�Z�ܦ�ޕL����*�G�T\C���j_g�D5|6�O�1b y�zO���s�f��T�N�8��9�*���S���8 �q~8<�r�-��_�	��bW�6ݵ�֚��`��?��eYԡy������w��[��7��έh����C:�U�8�,rU��9�%��B�`b<����:�wt�,�;��p.>�
by]i�B%�)/y�
�ƭI^y�kC�7G�~l�+��"�Kz�A�?��o��I/5x4����;��h~��3k�܆�����O8A��)2L��[]��*WH�8�9��b�w}�XlxVHYEB    2b39     b10�`w/�|i^���ь�}����m�G�����e�Ieu�M���b`�j2��9�g��5g��l�E�s��$!��$goT������E�i��.o^��PC�I2d�ؒ?_(Dj 1(ϵ�+�IOѳ��5��N���#+����	���JʆH�}�V�<ݪW��.8ꔆ]����0b�vQ4�1���C�ą������J�%�z
�����Kk�ؤi�6�x\�f�����|}�A)�[�M><&�f�dK��� f�^>a{��majQu8�aI�!��2�dQa
�o�2���Jr|���X�����jۍ~3bǢ+�DR#��Y.\�w"�;�hɻIf����
���e �k�e�v�������6ӟv�2��\��6hu��� ��0X�����YyF��*����u�=�r�\���y|�E�^_��Jɮ�4��
��;�H��)v:-���٫�'�$�L�6�t|���k�­�h��B�7��=�w��4���Y8F]�� �bT��-E�O�*ؑ�0.|2&�j$r���:_�4��V���?���ƏO#1u����Ae��s?�4�w����[-�5 e�\�/t�� ,VX���:�py��`F����QLk� ���<ΓA�:��}���Ly\!� �toZNȾx,_�U�WX�*�h�t�ԭ��q �t-�76�,o�/�1f�0��.�lA�XdNW�q�=Kx��O��}Sf�o/�O���s(�b�#8!4a�y��s�̼9�}�~Ҡ��0a�β������S�jTzS�������q��~���.�6����XmeS�'iM-���*}%�) ,��k��4��u��9x�;L#��n��::Ze�r��إTX��̔
�M��#�������
�ț��t$n�i��`�s���N�'caau��M@#&-���Oǲ��D,9�� .�ރ�Z{7u��z��D�?�}�<2��%�>w>z�Z<�i��X����Bp��=���d��m��>�[���:~�&-ߔ(CU��X Z)�q���]�!������ ~�:�>Ǆ��:^���Y�]x�yq�u�s����y�C7��D��;�`����+��#�pr^T�HQ�F�5�_�2&|���h�l���툧C�&�$���F�q���芓�o�d��#م6Z�Xi+�-U�;��$B�cr���@`�֧~�G�jje#�=�����~�Ñ)�R�a�p��u�"��i[o~�������$�h�}��~��l1�aMA=�!�dSJBP�y�  �����Q䊘�%x��e	���F1�1#̛�� 2򙛺�r?�MZEj��w���o�O�x1AO�!���m7x�L�+w��(ἳz��x\������-��=��э����F�� ���O-�j��F��x�X�]�������˔�~V��t9c��G!�Za'���{ʍ�z�kO�?�1)�G���793KoaN�pB�l$�5撹jؿ�@]���d�4�)�-9��j�~5IT���� ���z)'H��UL$��}j8N�[o�"9>k#�y
gPJ$�TK �p���
or�E�m�`D3Ĥ���M���a�䓟1�(o=�R�N 
v�<�_�S1���wҼۤ��cQ
]�XU�`�ꏌ�Ry��<��Z�د4��]�"	C�򵚋x��%����S�0�?�'{���卢����J�X}��+r����ި�iqw�+�M�
�u�I<n��1��|�AqM�∘�M��~�a�j��Ⱥ���x�|@�՞[i�[|r�#����)��]��ה�"��1�9�21Yf�;�5}���g~�ߚ�&�]���XN�/��'�������Gc��V��'TEZ�\��Z�"r�$�e)s�Q~��8'=]�s1Ǒ��*8�AP,D��C9Y�PzCHO)���t�_-	s�o4�a@�����69�?�Ӊ\+��b �NU{�jl�q;tcB�-�Ry�u��9��:>H�dR�	��{]���\�3s��|T�_S=��q0�G�N��}�#0�B��S��#C���B^X"ej ���=�����ճ+��7\�H�%�
��noï-����y�C_}1��o���^�@��TH���|�-mer}�R����&��aS�ͤ@=\���T3����`�S�4̮�	�����Pri`��a6��N5����WB\+�s�a�M��n`� �H`�S�{��SU��ѭ�����������b����úaŗ$8C��}d�_��C(���^����--f�������a�FNS�%�S�VV��0�kpr;��H��{#/
��I�q�rR��싯(��]�+>�S����MJ�		ۼ<j��Mism<z	pD�e�o;g$��ŧ���c��U��GJ��:������j�/�g���b�N�� sv9�9��õ!��A6�OT����m�0�����:3��S�[�t)~�ٷ#ƍ����TJ�V��h)7�� |��:_˂qc������:�d�G���\��"��@���ޗ��D8�%���/�9�OȐX=��&����6�Ov�#�dE!v�ʵ{�mqȯ �Ua���/�@,��P�Zz��$&��Z=r�s��������/�d�"2L��,\6�(�3H}��y�z�X>J��(�p��:=;|1�N`���ɿ�n�`�F���1�.9����YBf�6���}%�[���U��T���*�.�ώ���Z8.�w�Î���#��b���