XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����69�H�9����.	:�{wo�N!5�S2�e_��ᄮh�U��͕ ���`��8��h����Ĉw-��4O�#e͊k��ɍ�R�.)�FO��!��������$PП_7�	�Va���p ֊7��̛�kd}�˅Z=
�d�Y�jWu��g�ߴ��f�ޢ�h�ZePL�5�֟[�L�c�Tck���fXțHs�uP��>4��I��<7�#d,kR���5����<�E�kiK	`����R|S��f���my�'���+�.��@��ɏ��c������� ap�"5to���� }���웆#���9K'���H��Pd"��-T�������Ư�	z*}�I �7p3�!���t�a�
��ȵ����tr[���j���>Rv��ʢ|~��Hh ���t*~��4�j���!������ٙ#��I�?}�0.�X-庺���?/Pz���!���Y����hq���E��W�2��5�� h<��J�s�b�,�$E78)���OU�{���v��䷚���a�s�v�dA�
�N���Q�|�9=�Ox�61ͮ~>��i�$����{�r�|�(o�M�	��l���sǾ�<;*2ȣ��E���"u�������~[�&Η�C�=^ �8� Ԗ}ȁmJ�E:�ڣ�__R�����<�h,�����yϗM`�җ�
cv����]l��h�b�nJ�/TF�,7x�f�#��H�(�M�AO�Q7"���B�UE�5�)9P�An��Q��]mXlxVHYEB    1959     920�3�-׏_�	��X:�Y����2P=��׎,��i�����P>�˲�;D��:� 	�B>��P��uo�:5S�_��xN�7#қ�D1�,_�j���W� />�KaԆ%�V�-�1� �7��aM 	xBn�����."B�E����O�^sz]Ph�].��G0c��A�'o�˩�$R]C�1�1���IF�Pp���O�p/������(�r��6m|�-C�ڬ��nU}��k�Ɇ	V%D���=i��#z����E?���3*�I)S�9���q|J� ������C6q���(=������}ZK&���G'��z���X�x�
�&@�(_0]�0D�X��m)�����~���}�z�wy�E��9���,�@�@'�lC��@\k�;p�q�ASB��s;�S�ἲ�����vnz� `!K�cR<BQ�*HN���c���a��l�tE? ij#�m��)U)F�*PӀő�q�D�>R�M�d
)*\��>[վ]��8�V����k]E@X�z���Ŭ{���('�E���Nq!�7�;/�n@�	�྘�����������0(LC7�y��qĀ~M[Q]T�XRl`keKHz��x᷀�eFH~P�3�����3�a;��S2�}�Cߓ�V1B�G]��&
&g��Ꚅ��V����Sc��h�l���hJY
r�S��ƾ�v��_��Ԛ����2:�z��YzrYܙ���~1|�{�zf�i�/X8�ƪAк�q���?�I]R�eN4����(���J�t�crB��&&ͧ�W�ӨϮA ������[�a�/��@��A�� U�Q��p��쌀��O��
C��ɧX���r�T�J=�q��賹�2� �,�#{�"���Ե���������]�_B��y���߭��:��C`
i����m1� ��Y���C�V��*�5Aǲ�3^����N$���{u�\��s�c�֝0�ڦW������c�����0��ު{N�ޭ�@8����I�rT.�% H6�A3@:	*NZ�Ė���o} i�5�'��< G�n�ꀑgؽ4>m�-��>`�_��-�oIݧ	���e�溣�y��!����-|7ۥ}�hS��21����K�$4�����č�����-h�o�Â�%�:�r����-u�>����jȫN��8ʆ����B��W��B(7� �#s�}c��ˆNu=IE����G��~d�t��̃���s�v,F�!^[뜻�N�Ǆ�q1���~kF�;1���4:?Ƴ�%����NM.qƊIh p�{� �?����ð��y�����t8�ȞѺI������Y�gP��:��_@�5;�7],6 H[�R�H-S�怍9<�'�0ĽLT{�$�^'�h��cr�+�S�����_����B��U��h�c\�a��LEx�G��v����A.$�G��p:Nu�@۹$�P��k�{32�5�zSt_�JN���#^�h�2T��7m��+�VgݔU	=T����L)1�<T�Oު�0f��1��R��q@ǅ�$�R2f�z̐ks�0Ck��eûF��]�U!��*΂F��L����HE�\�D�=\qY[�G:2F�2�(�GU�e��Gz	XF��	��t�ǋAy5�E�j��a�=K���Td'ǀ�ن�ռ��ݺ�b�BҐ��N� �0�f��M�.v���l�����F��N�n^%ִ��%-��j��অz�]�B#3�\;@e�Z�6�Q�v�s�+����T�Wk�#G���F0J�V���*���&�)?��!�J�y��ѹ˸�A����?��>�o����*h�ܮ\gUֻB��`A��5�ZZ������L�Jm)�G�k���qeRե#��+��I4�r���Z���T2�d׹X�E?^�3f�@��cg}�n��RPպ^�?	�>:��}��7]�H;&쫻E A��f��oD�u�#ƞ�K��s0ž_���e�sݠ�z�F�Y�G\�Ϣ�cהF�Ñ��ˎY��o�F�U#40&6�"4�6V���5�ME�j��2�hy��>5>Iƺ~�%�������sETG���eE�f�y|T>��圾:X:PG<�㔄*1�D�Ƃl	":�SY�o��`�y��t��5�>���`(	r'$�<�ԖNp֪�}����PJҫH�G����	4�d4)���8*����SS�l@�����w�'��j�禲�{ � 
��PF���خ��d�[V��?01{���+W1��Z��@Y��op�J��NE���4��߁�|��Y+�eo�