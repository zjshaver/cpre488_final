XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��	��K���k؏�9��Ӱ.�݋ǖ�!�������˧�ؑ�o�з��a>��ۃ�ǫi7�c]��xhe����N��m���}k���W�2���\�Y[c�4�b�b'=)>�$߆��5o�L�An>n0i�_~�/>�3�q���u�'�yD�
i��-��?�2��R��/�D��JI�:���0�9kؙ��b���j�[�$������ĮPƻ�>E�-8A)�+�l)H]/�p�zH���Q�f�xr���oj��<��E���RUڅj=9Zs�����F������+��^$�������6+�+��>}Eg뺮}���W����!4��3]Q*��11T�3?^����"�V��a��dV���FD��V�1�Y�&k�2�#��{'��nR�؋6?{��u�kۥ	|��.C�� s�A��]f2e��7Lz�tR��G�l?5�-��+�����i��k ���t�i=�j˸�vJP$c2�v�s�Y~��)��&8(^�n��~��R�/t`c6����?Bw-��O���B���?FE���o�g�~=.�}>�\'�D�J0�ú�JM�.���{�K�?��Ng��s4��؏��{9��
�D��9[��+�c�i�'cfr��{���Zw�~91��x���ĄЖ��Mj���V
�G�d�t�Qn0�w��1h���7� 7`��[7�1o�@Cm{Bv��6qm��_d���7�J�3b�Jٵ���y`Y�1��Q����U�XlxVHYEB    374e     ea0�3��V�l=M��C�����d�Yu�ۭ��_a��]acȀm-�e\�`�mj�ņ1[�)�՜�y�2y�"�ƪ~�Xm��D̅?o�F���N�D�cl)0���h�pOU�F1*�M�T��g	l�Jlf��'W�4X�9��w� �>�}�M@�bHM�O��jU~nOԧ&��8 ���Ӂ�pH�j.� Ĩ���ȤN�����ҏ�ئJ�̙"�����֢�����0'�D/��]��nqz
	�v�s�B�hbd����`��h���a���މ�0D]2@t<��:�G����0�;$f�!ۖ#��C趂�tb�2P~�ޏ���� �UV�s���XHú���By�gL}��Y���ԗ����s�r�/�Pn�r��J��u�Q{DN`�z�:nA�@D�B\��C|��g
�Q���3�'��~rQ`.)p"�ƩG�E˹؝~@=��NL���;Q8q����=Z�=�J���0�-�h�j8�i��PGS����gZ�@���2��d�\E#�b�S-���	<qܥ�b!V���瓩�$�䦵(�N,��������z5#h��du�f�|-��g�rjI�=�o/9t��4E�3Hj\vW���!��,����=�8�}q@���S/�?��F ��$g!�Mi�\WI�A[��*<�M]n�ŗ�������)�k��`��4�M�����lP�Y83�zVʖ�V�`�fj�;�#��^��0��g�O�U�pVd�`ʞ��P�P����̉��#��QE�+q���,PG�gr�o��dh����|�kh�L��(��^pA�a�gŪU
V'f�w�ܢO�,��0^�ߔqٵ-�j-�����̜0H����lQ�=��`��*� S6�����w��� 1b�F��M��S��c\��j <�b��yx�Ih��)E\��e+c��s}�R1z��c�p�B_�F_�nq�F��p���P�a�Fh� �@�k���p�Kn�S���մ��d.�M���	�B����A@�
M�H�r��z�C`�a%+eA��E�"D�[�=!v<�G��i��C�o��}��J�(
ɴ��(Y�F��ϻϙq}��s�� "�(FFG�*��ͺь3P?x�h��9x[A��sZ�����2T���8�'4��İUcg�\@h�a�ݾC�mӅ�B�@�2�	��zg�.0��O��͟����ޱ\�.��F�Ԙ�J��e����Hͣ�7p`f���2�5��L�����h�r���є���ӨK��-}�$p��T�1"�2��F���K ��Bdp���w��dZAg"\@pP~ȹ\վj�\UH�5��ZbB�M21�󾿈D����y�_�Uo����
�C�d���A�:�f߽��@�M2���R��"r1F�~W	����-�Gn��X������ґ������m��\�
˛�j5[Q�.=�+�8޷׈̊�݃�+��� �|'���d����<����&X�N��B���9;�hܢ�l	U7�6�=ةJ7�����y_��2PT3�Ec��%��P�BD�E$`>[�%o�����֪$�l|%��|Ot�����C�����lo����H�K�� _�}[��s�p��?bE5ڢ��j|����h;^�`�����P@����bg�_���p�e���8�����2�GHR��q�Rʓ�ZP�e��p�fZ�b��6�O������܋�pU��l�x}24�?]q+����Xb�ʠ��CSW�$�.�L� ���$}�����i;S�����V$
si/�׈�mz�6���UcR�p6�;�] @��Ƨ�o�</��@H�f��uX�&W�VhW�t�z����_'� 5;��ډq2!�4L�PJ�Oi|� BU�~�Lm�q}I��C'�/5/<�	����p��M(���6PW��23Ai
4\�ʀ.��-W'}�)["�o�"@r$���Q|ݮ�N�4}��U!)ʳ�_o�ʻ�{W��4�De���g}��4i	�����̦�˃��&���|�{/X�1����&��i�=��3;��L�>i�O{3�,INo _�������9ڂ7���@2^��;�	5\	�.�|~�p�m�/�91k�v٪�j��7Uʍ~�3QB��15m�H����������BW��s��4qN��!��qbƹ�=�dn�e���06��)����}������ۿ��$�ff�w�s��M��+y )#��ac�+ye��c�r�72�\e[ڏZ�ly�r}��l���B$�8���1P:e��Ż�N�k�SK�"!��w_��$	#W0����� v$7T��� ����I ���ƥ_4i�ZYW^)�$���(J�Ѷ�.��0\ K�p&�&�����Tk�֘�N7�t>��S��vY�#�����S}zu��H|�Iq9?�lZ�*�nH��ٝ`F��î�˴c[��T&�M޷�U������a@�>4b*Z�D�2�����3}��U�d�Vŏo����%�F��d��_��b�M'�2 n�=D�l�f�[�]�Vۓ<�0�I�nL;�j��V� &F��`�O��(B�	������q��
���x�d�-[����.g�"I�`��g�jmku��eJ�ޑ�Mi�����|%�Yj`��z=�遄8{�}���r1�vc�*�~˛	��E�H�:_�.Q�$hB��E��#�{T���5i�F�������o2�>$����.X֤�&+�p=Un�1�(�����u�������+6�Ȣ�v�lD�M	��k]�� ���Or�B-�\�27�懄�����ŐX��G�8f�4B�x!��_������0_AvY� l����=<9�ήI�r�e��B���S�L��zO�rkVز3,3��zm&�U�3� ���C6x/�{�� 壎��\��5-��qyT�K�[v�gD>�谾 �/�@V�%i��Z;��O)���c�ȿ�J��M��ӗ*ˤ���Z[�]��2n�2#?]D� ��D�f����YEe��(<��Tu��5��#xo�h����mj1�_��k�n�V��V�fY�
�'���Cd�G����[� ߦa�H�g�5�t+��P>h7���l�+�U�����V]��An
����!<���Լh�#�����u��4����;tm~�,��{���v=-;� �~��#u�wDk���w@�6�Y�(�'��YFF, !�Y���ث&Q�+Fw�;
��%Z����~�x-Z�d�_]�Bn.wyT���J��Ż��q�5 |���7�u��HJ@	9C��A��	��Y�����������+�Pl"�I���P~PV:��%hR�c�2�;�V?UZ�ʜ�S����k+��~R[x���@���y�̲����i2q�5%Ie8Z˂��~8���n�um̀��Q� εOܥ��zC�}rtBx[ɭP��`y�-_u?��N����%�o�JxWZ
-�&,��tY��Uֳ���.G�_��DB��'��R����ǁM��^�U�@��G�Ԝ��Q��j���� ���E2��]J�Y�+��x9'0�����x\��0p}7X�N��%	緻����ֈW
��m���t�����
My�#z#Rn�*�����'�$��9Wk�?���S���by���	�9���|��b \���