XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���D�5/G2�ifh�A���
bǐ6H�K2R�+BN�t�v�^�5N�������|*���O<p�A��Opf?���&�T��h#�s�F{~��Q��3���&�l��p֜b�"��TH���YM��d�Q�hdN�<��M��ß��AW��<��H�)S��7ѽ�����B.z�RC'e�=-��:�s��9�~���E�Q�r=tv���Nɲ������Rs�_z�
|�:k���--�<.��]�W6;�L�O4j��3SD��Č'�L���02��ݼ�O�ձ?����0[�%���Ԕ5�,�����H[��!
�Aw�����`�T~r{���S��*&�S*_��Ud��5X:�kⱷ�i��P������:hf��k��x�ʨ��ϰ�;�|�sTJ-������H��y� ��Sa�V}珈���H���#�1�<_Sv�y��	�C�R|���'���ٸ����(2ۦ<C=�=(�M�w|\޵p+�*>��Ó�H�g�w�c�*n=	'.{I ��D�����y���/�	��Q�����]�����9Z��"��H �W&g���Ҡ��5-�`�"��h��R�%I��1f��ҩ	<&��=��MT;����],�]�&8�B%}v�<�hl\'`6E�Q�|gNC�x�	�ڇ�ۘ��ΞL^sPw�
"��1����������NX�v?�'�kP<cQWțǁB��^�F��V�o�#���þx ��1S����v�XlxVHYEB    76a7    17c0��>�P� rg��N���w$�(%Kp���e4��x&�Xu���'j��}^5�fH&Z!�s��J��od: �*x�4��z���L謬�?�����I�������X���L��:u�!Nΐ���%g��p������)�%�,(�`H��QH�w�8c�����[����y\����xG���Ŷ�_Ie�߃7	����-�=��7D`DN�Oy� -�|�(�
�D_��}=:�7��H��.I��L�*��%��r����$Q���}yJ�[)���{�m��E�#��R��f�Cŵ�<~��@i�4*����Y:�@����15��Q�Ga0�sy�׋��ӷ�Lڀ@���Ō�s�v�-#�Կ�:�k����2z1�O\w�f��m��&��/�ʝ����;��W$�s��~W��X�d��B�s:t��ܝ���D���y��[c����{�����[�����&�OHC�k��
},A�@��UK��&dĢ2�{�a��B��d�����G@nt��к�s�j�FlI��h�dH`R�������X�߇x.�5��ِ���,p)��°�T��7a���6��v��jŮ���8��M@�H"3&���0}�|c�I�Og���]|�4����C��	=F�l��vy�zݤ	:'�U�H&�̛���o�̴�Z�y��k�R� �b����Oƚ��S����6.�Ș{,�A({/�v��w׹Hf�ǀM��I�Ƥ��l�Õ�e2��8n��U>̹|��v}jA�DwY�.Ё󶖵�#�&�: t_4fHk��x�B,���g�7��^����
]�hR�0/~`�I���h+�c����L��C��Q�V�6�jN��2�3�:�	�	�]D��4e�������zqu�D�ro[�Wi�������v�E��Ư$՝х_7o�u֔����r򌥸2�rtEӼ�Ƴ�GE;�[ͅR�	]I��v�i���X|X���T�w�]��|�h�d=�����T��v켵�D;P|)ՆD#14>H޲�mvI��
 �}:<�G	��p��-t(s��v�Ў�q�U�WI�z4�nL���@���D��U4ޘ�=}B/ˉ<��ܼb��羂��I�K-�����4�@>��i��߹5J<����?�|�;ՔuIl��'w�ZT���s(=:��QD�������AM�n����B䙧�9���@�Ϡ̱K���/i�^Z%v@��g�;��~~�Ҥ�p����:�����������*�F��?x�W �7M7蔡�F��}���"h��@$��쥆��K=8��S�IJ�H�w2X}nt�~0��5\C@Z�_�z�	Aq��|E���9���kF{�`tf�#����s�M>lc�~%�NaY��t/�;�:
����	��k}pn����4@C&��'c��IWUS�
@�*���Sr����d�mL�� �ZU��#Bz�}�B�t���7c���4�Xe��)��0���#���^d(б�ݟx�;|jx����D�UJ�����(7-���ɇfXb=�@�x���MNF-=���Q�Sx]/be]���d�@l7��J�	��z�yȈ����q���v�J�ъ�_O���R���Y��0���҆���_�Rk�&f�,"����^��;�׫�D��u\q���N	X؎D�~����*�����Է�iZp��
��c�7��x�:���e0-����[��|���me����i����Y�]f/�?������i�g
?�G��O����.��Y s����E����aT}���L�p:�k�3:���'؏�m.��t�9e �-��7WH�H���TMw�ʞ�TF�*�8�����$�pK�(���;O�����XQ��u��5u��&��6 ���>�lQ0��#6���8���]~eba�����6X��J��h��q+��G8�7��:7��v�Ќ�5���y,�&�{O�:�p�hl�Oh���*���m`����MLۈ�+��S���f&��
�l�K�������"k�Z�[V���҈�J���Ƕ�$��-��[zB4��b���>�e��?(;4��-O���%f>k�6O���T9��T=<����Ky������X�����󼶾b��rTJ���3�Sf�Zi��j�������?��?�2�@6�r���5��\F{%e:�۷�V�D2�F'���yĳ]̼�;@��&�-�MҸ!ߺ���"���W�F��K�҇m�Ъ�yz,�N_�[4�X��Հ�'��Ԟ1��u&���W>�|���'f7�6t;,
��ڟvK�_+U@ ��.!rD��E/ ����C\gݹ�r�x9��
S?�&��%�����UV���O�ŀ#��㎸R�;�_q�r�~v=���h3�F���eK������@&{"��m���F�A0�t��Z���:��M�+d�.9�ag�<N\&Ű"^��Q֕��(TL�P	5�`o/�U����ΰ�(\��~���c��9O�#��C�*�o�,������9\xd��7���
f����f��e�N���!��^6�Z)`�� 9m�`���r,�ws� 2�~3��zF�T��q���5@��I;���@A!H��U[5j�T�ǽX�vsQ*.,7��$�����j˦���� ��퐇�&1�#"��vW{��ۓ~��ɸȘJ��<q��^�2bK+�L���v����_��c���^�t��`f�S,R���s�i�Vk�C�\�hD�+��3�|�&�R.
u��‟���]l���r%�����L���:[�d�~g���]�	}��
�xcm�P���Zw8��F��;MS��W���0O��}F�a�.��N�;�N�t�S,�sh��a:��t�I��~�ݛ�3?�Ap;̡5�s%Q1���^�K�+|m�ɹ�f$�/�>�fM�sY���q)�(����0�Y��F�Q�={�0�W�X�tZ�����3�I����kУI�C#�����8�,���DV�� ��?']��ŢWG!a��e�����K�ÿ�����$��"���@j���^����5��⒢����#Qa7pS���&.JA+"�e��|"�䙑nدY�oM>3��.<�*�\6�uaTuLK���Iz�{HE^���QR�bV��x�7��QnM�͕�Z�wuGtxAc�ƄLOo ����_ŭ�o���O(�J"�'Jp����넯�D�҉[��q�(�&rǊZU={��{�8&�{"����ښy�q�/RC��q��t��#�Y��ć��|�R�md��U;����Nv%8n�������ZQ[lYNl��j|���)����qι����ˇ������+�L��ͻ�n1��H��Ʊ���Owe0hiK׍Ge����d_���>�~�o�v�)��NW����=��J�1J�W�}���(���Kt}�/M�X>�.R�@�5c�!�3��?z���a���������Zww�6����X�i����jg�j�h���X=$��	�	��ק=���->��+��&	�^���OM�7v�ja?On�υ_)���I�ٝ�{��+�TEtMK���Bq�6A�^y�2ۖ����O�
r|��;C
�N����P� 8�uC̗�Tk>G)eS"1u��&s3	���	�����$�`Y��_?uX���ڲ�k隺jɶy1/Sӕ��/%&ֆ�	+>���Ɩ��H�v�i�o����7�P�0�����_v`޴�Ȓ���u9��:�N��	�Q��ZIiUVB�Lm�'=��;L���oU����=H��¾w��L��ˍ3�}��n\��<f�r�׵<1"�EF^���E����������_j�gN[��U���`�a�/�F���v�F��o���~%M��,Ǿ|�.}�J�N@o�pL�ҟ�JDUƴ��px�`H�7�?W��;�(	�� �̫v*~?|ƥC�����X� ��%�堖1`�K�ó\����!f���JSԁ����>��{�	����S��2U�̇d�_���=������I�I2l�{G�WE����Q���n��I.U�t�75��Ѕ���Vc��,�Mk��͝Ep�H�� p�c5`�[e�:V��`���
�����CqiF�i"�Wp��`��Q`�c���$���anv����qI��F��(E}i�6}U�9"�r�ņ��%>c4����������Bۻ6D���\\I���Tޙ��ẐR�9���$�E�ˊ��#2?2*g@@9��a=VhK��>�*_�nR�� �J�Q4S�����Q���%��\�v��XV������j�!��APT��H$��XW�q���'��l6<�.�!�C���[f.��Ӝi�KG��O��x�qF����:�,�Z!���s|��(ܣH�<�+m�U��]�l&V*$��f�ߛQ��S��ޤ.����s��=�<�o���/!�A4T!�ؿ!+<X۽w/�sG���.���1����k3��^ޫ�����H6�[���yoTC�s�㑚��hS5
�p�P�
V���"��E�fB���2T\�P�D���k�pY�,���[6F��.SHq��2�r!g�_��<�9�%hi37%[�"�q�Y{�7��Ɏ��w��^pV�)�O�٠�W��ݡ�6��H5�Ș���A=�๓r�/�v�|���P��a�+l���L�MX'm�$�-��H_}Uw�Փ�`��
{��[�������@W�aD�cbZPl��.��P���e�ݹ��'?�ڔ-N?4{�x������_Q;f�0i|p��I�ϫ3��AA�fG�d��VkQO-�_�p~��p$�F�;�>j�m�{���窠�&�����a�V��Sѳ���C������^�Eip�'k���4h$2z�E��?���g��Bu�^;��D��/9Q&�TcУ�����y�l�`Z�ĉFY}k���N��l�zcO��-���jW�����ݚ�P03{�v^qS�x��ȵF(Jba�i0~� �����H�p6�z���a¢4�6���l'CB�����4���O+!X�n�����I̟��qˤR��hs;�����t���\4�]��f�NJ��\�V�4ifb&x�s��iܙ���H1o�D?l����|���"���x����I���޼J�mi]tɦ��HhT��;P�!�Y������ �\JB�'0�����XPz�Em<�t�Yդ���%*uZ���Z.瞋�k"�`|ф�r1��Fu��u��n�S��S_�%π� ~W����3S/��c�����Pp�-�q~u�۪�Z�I
\Mί߉s�Zӱ=ZM"��|�N����y!/����~
ɢ3uS��Py�\�ˍ��gG���^��9�N�ʡ��P���� ja	TwV�u�]���ڠ*|��C����b�+�E^g����?���+��B/Y�����!x����ȗ&�^���}T��k@��DA�0%�6�N�����9~�k�3P��[O��Y���"��Q�0V|��8���}�.�	G1P1�گ4��t��A1WP���jToI�['&��ւ�Ve�Du9�����T�2�����_��#W�1{I�G=����.��ٟl�AL��0����x`r�e���B�w��M�h3;�*��F�f�+����/J�1�)�9�o,��yAY��a���?P�ؓ�j�<�ѫ#+j NQt&Ґx}����ޤ�����{�����:5���P��i�&���X���8lG��g���������^Vl�~^���Uw�,F@a	֜���-:��w��%�}���<��U^������,�0K���������o����)�������N��m�£Y(M�Xo���F�q��[r�ş�ڛ''���(�n�_�׷,cBؐ���(l�P��ڇ���O���Q��A?�:lT��V���=�Z�N��K�p�^uׄ�