XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��)1�
�4��h�|�k����l�򿔯㴲|��QC�������P�S���k��%��QAj:�"S)�#|İ�E| ��8�Y��������	W1"����K:B!�o�xg"~�':�+A�C��B|���H��%�U�5��&������0@�|}���#���RB%��B�&��|�T����r��=�C�����z�����̇�D��Q"�,�,���|�Kf�� /j��S{���+�%F^VpJ詹mITϙޭ��4 ������]��:�w���9��.�h���k \��4?���Ńu1�o ׂ�z��.�Cu+������C$.��o��<?��
���3��F�?�~X/���:����%�EӖ+1�b�>�W�x��>]���d)m5��\�:рU���W	�AmB)u;��xf����+���41���Hd��L�E�u��Z �G<��<��:2���A�X�����a+�q|�|d���~L��):�����e�A�����n�	��Fx��!Ɓ���WRm�7��&b�G4P�s�6;d�fw�b�U2ؠ=@%a�dQ����H'�<���R�M�(�ꉥ�oq�~KM��_�%N<#�G�*��]�k"�+��Wʃz)ӌl��S�<*{��eHp&�ܑM�����#J�tS~�0�g�A�]�NlΖ�N��~z�+4�'���'�߁���]�*�Zta���$��6+�-fng�X�-y	��4�֕��p6*/��4�ߏx����/��
�F9ql�9��_Q�gXlxVHYEB    5d54    14e0��7����8�Ǹ֭�;`�K�Ò���v�mDoW{�?�m���[�L��B�g��w�m8fZ=�d�?��3���o�V�s�y_�����g��z&)(�Y��՟|n�zM����Hpy�n��?O�����r��yjK �[No]u|�G��$ ��>t�N����TH!%��϶.�^c/9 ��8+��%I������D����r#���۟�^[L�<�8��D>��Y�-!�v�lp���2!����Ah%�%�Ώq@�1B��ԉK�i"D�G�'7#V�K[0Lb+���)���e|��Z8�w���/z⦼���[SMeM��H�q�����2,�p���m�:$���C�3Q`:I��̄�����@IQ��<�_��)�Ծs�i�C1�UR��i%�D���]w��'�!%ݹ��FƯ$���[�氳�g^�_�CA�U7&�f��u�����T4�NT����_�D7��[c r���L�t�I�!V�#.�M"�����8W""f�ܺx#h��C����{܎��+��}] /튄!��a�� z}�!55�
�Ĥ������`��D�<�̢Mjck�F�L����5c�h��S?ߎ䞺�i��%�8�O/	�����Rg�z�5��[�x��O;1�Y�*���? �J��Y�_K��6sGT��%��q�t�����J�@z`�	�|����Е���D&�)vD��(!����7I�i����-��W⽘����~s�Hoۀ�_��B�-����Mp��+��h�n��I��׸`E4�f��:��d �	���6u7� gk��uu��׏���������CV���Y2���oy���A!4Yk|a^��¢p:�I$?���4`H� t�������1zp���T`:'錚�g���\I��:p�z���f����j�Ҿ� ���g�Q6��*'�E"@�/�����s�S�NE=	s��;L���y]�$S]���gX;+ ��xGvА���4��(�����l_)�fЌN% �_��-3ߙ���w'��]e��ʩ�5K��$>���ˬ��;9|��_)��<�l~�
�;����>���3rE\�P����5�/��7��}�r[C�j� ����j��d�(p��&������3�([�ՆDB���	p3Tv�>r���\�άk�z��4�j�(��mi"r#-K��]��>he/#�e�~"Ƶ�Ym�[�/ٰ�Jײ@��p4)V�J���B� C�q�t:�p>Tk:S��(#$��Zr��+�JV�nW��f덒���PL���s�o�Ѳ*����Ł�1��́�&��jž�"X9��x*T4fG�R'єppu�3M=z��r����0�u��HY墩�:�|>�/�,�7�#-�� kV4�۰���?t˂7�0yd�����������鎥�2=��"g)]�>=@=*��;���i��B�c}4�+>�H����
�!�׸�������](Ze9U*����A�3t�䒨���J�>ZVS�:ǵ��v箯��7^�K±��Ҟ�8�%�)��נ�Oc�g*iu�P�1���.7V�+rh_�Y��B���Fȑ��s�P��,��S]���ϔ�tB1e��O��<�%~���n��e��.�k/����s�y���H=E�M*��%�������Ʒ�B_%8��$}JQ=��D�U���^�J�`p���a�"�6�vM�������S|9Ȅ���_�^f��H"� ��-H��Cm^�����q%���Gu`0 �n�wp�u!��bx;��wut6�3���g��P�6G�����^{�k���cSҴﱞƓ�ϷU�]&GVQ�U1z�gI��k'�S6~W�Ghsm��Z>_A����!2��x �0��\<Ý�����r�U���]��1�H3�l`\�G`����2P��S�d��L���μ*wWzG�oՃ��ZΫA�U����s)DB2��86�j��o�x��������k�Y�>���\��i��eu��]qS]���eY��[�C�N�<��(�{*1�i����1�v*d���n�|��P���@�t�O>���#��5����a1�2������r}�ݳ���`[��vx�h�0R;Z�@B�>cr�q���O���6�s�Xaξ�B���l��cZ�WY�)	����X�Y�e��5��w�."|5k%l�b�{�	�����<����b�\��-��t��@8.x-��M��v����&��򼷇C�d�ڂ�"'��6΍ԤN*L	G���W'G=a��Q�2w�����@X����oGYi7m��!��M���v.)t}�27�yA��[v����@�F�D̨#J�%p�������,E+:�Z~}{�6B���9�x��{֯i�0M@!J6�J̌�)���a|��<� �j�j��M�oG5&����$MgSwy��K�~o5:�61s�a:} ��A�>�ؼV0�^VF9�$B��w(��8M�`dB��4�����߄[ox��8�n�ė�|�lY򏛂"�����+*]*�UN�-&bՌsl�~t�z��[F߲�'6�����$e�p;?#K8�,'=	�wNY��?Z�YL0��Ok ��:� ��/z��%G[�q�����,9$AI�P���4F<ҠV{�%�f���8��8�艄瓷��>��&}�m��3��fD�Ey�[�N�`��f6�3�O��o���CE��޶s�3VȆ�uv���ZSb��|F;mR�HcG�<h�
N{����02����g?U�p�Á��'�Y��͜�|w�=-�<�����H��٠b�~֬⼧M�+�D9n�QX�3�^�F߳�k�e0b��G�e�E|u�{�p^ľ yі��1�P�	���Ǟ�E(�r\����� .A�)��L�H�q1���P�b�z���-SĬG3��<��od���Kq+��x�%N8=@��=%ʼx
�i<�X��v�V�o�d��b�yoY������Q����]����Um�j��=JFA�a��`��᧥�[đF�۞�^w��pC93ZJ��@Ts�ѷƙ���T�>��R�* ����-&���a�����&Q���%�k��F�J<U��6��V ��<ݲ���UR.f�Z 0ZZ�݌ $�*�B%\�ϱb���,�H4��LK.i�x�= ���y����K�L@�Ga%�O
C&�0w�.�5�Kv_;�Z(��Ŋ���T��[�;L�hh�,ǌ�ؽ�\��El� J">܊��*K$��he7�������#�&�4��ؼt4�-�*u�s�ӆ��i	�U^�~����0$_��܁gX$w"O���.��8_�T�����p���a-]���_ʹo�t�-�� m�#��ފ[���S�]�0<���gIἰ021x���O�gD��C�#�¾�$D����:.n�B��W����Q�7�NMB�{�ĕS�M��Gn:m�� K�x�wY6mߨGg��TG��~� _�F�j��6kR���nn!9�E&�����t����hK��A�M*]��������l�������_��������i��`�
����V��:�}\J�,	k\����b&'DE_I ��`z��Ԧ���[ �����bI੿s+�M�z�g�[��+�}��9�2nB��!�沁Bj�iuM�p��Zw)ٺv�8.<Hb���3NL��y���_���'=5Z0�Q��vf6gì��ޯ�*N����ת�.EYV5\x!�h���%��D�>��*t��@�5�o�����8��L�>Q]_�{2�
O6��O�����S��\\;t���\�k�~�׉m��9�YQ���_���E0�ʹ��7ώ�!���v	JZF�[8C|}p��g�Z�X�O��,����pw �,�����̝>�*n�F�U���Q5�=�0�ű�q����^������?֐x?X�FaS��N����^ ��ӗ�5�5��Z�8ð8�v��.������rN �b68&\c�{��Xp�ʢ����2���+�t(j+B �?��8
M�U =,oD�d83ʛ$��1�I�4�X`+AAz�R��Q#����۾�������@(���|���,X���W|U���K�B�t�/�Ӈ	ێ��=��{�N���{�q-ȟ&4f4���`Dݦ)��z<ց�k�p������ F���Z��TZ��Bbnu1�,��q�_��{n2�T[�С_ei�>��=�):�S�v�p���ߍ�5(.~��?�U��<�mv��>h�a	Tܦ{/��[g�4�0j��D�Y�� *�����$q0�ӌ��A��M���o�[�3�8m��oŨс�Q]�Ȯ�ݛ�WC�C�y�;A7 q�^Q��VP�]�K�n���\]��G�H\���|�ɝ'�����/���%���M�8�7�E����)K�!M!����F�ԻS@��"�e
�&#���/��p=3�+KQ��U���V?�a�zi�ǘMoqE�/�"mO��NY��h�q�Պ��jw����4���F�ћ�m����r�_�Ӊ���p�=܁��"n�$3/�E�ɡ�_�ꯟ'�%�y#7� ��J�n�:e���p�Agsf��_��^��[��зo0 n�y�M�}șH�h¬p��_9�ܠ���xW]�G��r��ld�l��Y8�4i
��Գ�g&V�f���P���
p�T��c��*"���337o�뉫��o���٘!���;����N@�6@r�-9�W�Q�3���?��<kećq���A/8Q]~Æ������b �_��	�0��}a�����bN2ӽ�uI����ۑ_��Z<iE�KG�x��Ю6G��am)�M����������7�單��ԘcS�[��YPo�L7�6j�4n� ���YZh�_����"��uix��%�bЛ�h�X	Zm�$��������kA2 (��.ˉ�P�ΔV��s��'Aթz��}�^��SvVu?è�D��NIK��s>���s�3!FA���c�2,�T��Gy�dJo�͟��|�K�)����J̉%]O$��Fr���J��An�|�o3�����dC�w�L�G�Z�y~����U��%ۊ;�"+j������v5ݏ�,�ĀFy�]���^�r�GT��l�Y�gs��#������s
+#�'���koa�+8�;�H������`�"�9o/��<�1Jə�����)��­~^�5��1rcJ�?�@�J���������xn���h3�yLH�F�Ԓ�ӧ��6���k�+����w�R