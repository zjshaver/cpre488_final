XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��@��RՊv�vi�vfKf����2�l�������r�O.���ݝ04��P��R����h>��7�,����eL#�fI�Ns/��f�0��A3�	�����3;��ε!k�/ M#c�e�վC�A	R��j ��zw���m���^�[����MG�]�b�f��?zW���~�)!Yp�~�R�
��q�&0F�f�����o`Ξ1�b���A[��cp���[kx]b��4q`09�cn�BK���P��G�d��s�fA(������Ҝ�%h�c�����v�+p�]�J��։=7�O"9�IY�&�u����d�&���%:Ù_ޟL��}c�zLZٷZ���ȠF��I�µT��N5^qis��ic/g~�8?�,�I�pB�l�Wp}�[q�R��gW)x�ψ"�`L��OΫ���s(����eC`E8�z���{%g$&B�~ߡF%)8Jf��^�X����1h���<�����s<9�T�&�]�ǂ�V�y�%��o��au3��*��&�7�8Q��2�lp�j`.��׸��r�J������Ru,y.b��j�9�Q��&��ϖ�.�ιO�0�Zh|HۆQ���U��LE�bVD����o��7�kI��z���bX�?�s��<�<���1�1o�N(�Ʉ}ԝ���G�V	��=����B�͎Q��A���cYNk��xդ���<���08���Û�/��>�^1�xa�1	��Ο��R�JS�Ʈ�����M9�J��6+XlxVHYEB    13ba     770�i��*����C���lΫT��I'X�����NrZ+����:�Ϳf߰��gm��(�'���7"���"�+{�;i&��@�4�RCM.����ߋ��H��Y�DZ����I���?ୣ'p3�^�ic���P�a^�����'r/OUktq/#���'[�^5���D�[(Yk�~_[��;7ق��Or��U�-��?@H�S�PDx(�+� D%2��g�)���:}�/"�vX_o�fRE߃ +���1����Ѷ�<�-L�ߓz���E���|l#��n�W�H�L�7!-i�3��*#�4�M��x@�TE}]O1o
"�l�['%� ��O.�����G��J�Y���E����EY�.�{I톔F(��_Q��x���^�I���}5��؝�_�)�� !f}ȡ�]����j��/az�K7�cÐ?����F��_�4�ʡaN��{����A=E�
g_%����`����v�*�����:��_��,���*��n��|d��0�\����9��P�1c��*3c�j���6�!A5H%ZDw);خ�璂����P�����k�!�˘[�C��(W�N�[�f�nGg�ux�u"7���f�1��I`�E�lEa�9��z9��%�Ζ4�Ԯ��F$����h�d����F�l�e��0����C�b���r�� fB_��ܳN�Ok�R�&�}M����X�� 	;�
VL�wW�A߃6�'��)A�yݧ]��V�k CZY%Q�q	�o�A��Ea�@{�I����Au�1��T�w�V4Q��24���J�Ԭ��Z��op!/��ʍ|(��/ϭ���QWT�ju?t!�P��7Q�����ZNS3P�@�`ZdL`ZBd��q9�wY���u��� ��#��Cp@sm�z�x?%��`�+T���(D��m�H?��N\pZ�'"��"�G�
g��|���u�;�:��U�׊�#��>f�Vc�q�.��ngbإH������_���$��2�@S/��ƵGk��Pp0UJRF$��O	�h#�w%8}�q��S0S����Ok����*��=\n8E����YY>�u��*Cb�8�B�����:۲��1[6��Ъ,bnn�m}���6^�Ǌ�/f�^�Gp�\�>��[��~�X�W��X5�^2��+��>�%����U?r���0�y!
8F*jM�A��N��+�poa�c�Y*L�+]�'x�����~$C	s��g.�Nh܋|5�`#�Dњ�[5����~-T���.q����i£�qG�h�b��NY�:W"9�de���\".c�BB��Jl���i�5 6=!�4��	���I��A����G\�����Sd��`J;�f��jϓ���O�*1-�&���*|�'UNjt
��=�W���,N�k������P� e�@���:��*4,,�̤�	��M�����Rpb�%2�K��˲O0���9���>���7�(ڛn5�2�>�9o�s��0�rW$�q�S�I�O�L{3n������������`�H&�}Z��0�v����^�a�S�h����SpYg����U�b�L�>���8�ї�KM�4}��K�@R>Z��O��i0�*�O�[�b&���
���F���;�3�J��C���X/�=���YbkW����3kƼeD�����_~J�/	�A�9�%���ǅ7��7>�i�� $����0�T�*�BD^�w_3.���}M�!��d>��'�BY�*r� �64��aՐ�6O�aF[N+��L�D8z�U<���5�|dq||b�[�����|�P���*A=���=�Ĭ���<�'��Z2����Qg9�YW@�$�!����F��t�]-P�v�w��<�
����Zʫ�՝PZ-d'�