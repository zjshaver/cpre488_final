XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#���2#��F�pA��L��i����K��ե$�nq7���^��h%���ى����( B7����o����>��n�H��oD��+5A��n@��� s��hx����C��w��^���n�ٹ���3,�+-��Uq��M�q���8�P��l�ӯJXލ�!����N�(*%�M���$qHR]���L�M������n-��+=��@@cy =�>D��鉐I�l\�L5 �Azs��j�:���[�2��Ta�I� %�;���*Tq)k���dZ��rZU�%���L���T'`�u�˒?D�q
�TFz"��W�z�������>r������7�:ߧ��6��չx��@ʮ��+U��I�xr��P�π}Z�-l\�G�*G�����m\[թ���iN���]�x��<`hH��S�o�- �Z-ˊ�7���\AD����Lپ���E�PWV���5b$���`��#��������� �e�5;Q��:���M�����O�Urv}��A��>�]�s�8�ю�tTZ9=N&���/JC �+�S'�I�Z��l���T��
AGs�D�h��3!v�{dzj�TF�|1Ն&���ΕZ��")Zo�©�^Ji��+l��s`5�e�3a�_O��E��Ϗio]g��̀���(�P5�%]����vSPi7��~� ,Ҹ���o��Ja@#+T���BG+�]�?��
�w�9a	X��4q�����±T�+Gf�XlxVHYEB    9fc7    1fd0ȍ����he�v}�����p�Vn�GPK�ް�m����9�XK�B��zA�Z�׾z��BO����e�T�:i'�߶o�A?��L�;���~4l}�V��h�����YNCz䅭��Qlz��v���a�/��Ntq�%�k~`5���n�u�����`~}��}������,���Cc�����E��=�Vk��8�����Ôᅲ_�v+r���{�t��[���t�93��}m�Fm��M�5��ƌ��4����y�"`p�\r�Ν
(f��&ʍ����l�s�3�t~�hao+�=���y�eXo�F�ܭK�U1S��.���v0�qW���T��,����b��*`J:�%��%����~����%3�&�#Q`������N ���>�ӁdB��J��'�Kt:�dx\�6���f_��<��c>a#��¶������7��8�6�c�C;snO�娹��7�)�B�!P(��R��i>=��T�S�0VM���܄vo$h м�@�e�j@}o5)b^�R@6�̸k��6C,��2\9RQ1�w�n*<�)�
Q��}f�U��/X�A�C)H�ĳ=�,���<���������j׶;�W����$`�T~ c�����Xs��Ig�CL�!�T�A�9xT���~��~��ش�k}ڦ"W�U*}�9�BE��	D�c�Fjs7�#��J,��$$Q��>J�ˁC�ɀ��Wr��5մ6������H��5[��������ϻJ�Jފ��ѷMm�Sutn�����p5e�;�}	��2�(xֲ̪���u��!wM�H"�3��'�12wK�&�G��E��U�V��f�� �;�|I��K�7�|�+��PHHIJRy2Cs4�Ix�FRws�E��9�dndEk�tyI�w5S֚�R�m��h!�=U�O
q�7���Ejs~,�ca��)��rěT~��D~�bۉ��"&�/`�l-9�7�)m�rM]�g"��GP�>�ej�W�R�S[��̯͇��czq�:��.��zl.�k PQ���x�R����m_;��X�O�ЍQpHI�Y���9)��A�r����,O�?^ANk�c��cE�W��%�\���V=^}�Q���	��3LK����*�\h�g�D��`f��R���ީrj#=���_���\�Psx��Xn�r0X�OM�,JW�.L���� Fip�^�����A�f6b�X��(C"b��&���e2��������CX��W)�O�6���u^=Ȑ�'r7�����*���l8ԙ�5��=f�m��Мxy����ڨ�T���8,@�z��h#ġQ�����3 �Q*�@u���h�k���:��8u�ְ�W�&W@����4"b�K�&�7�����퉲m�_�&��j���S%y�"�+Ŀ�o��!�|`������xq]��a����TMk#�g�~s\^�L (^ $Ǩ��l+]�U_~�8c�#��
�CSQ=���qX��9�QA/.T	Ѱj�L�cT1��A�Ό��i.S1�5SW�
m�7�Pq �n�TR�"� �!���Hxe��π���;s��䧙�Y{oG҉�V�徹�h�Ih���K&���t��"����m�(�_TB�E��"E-�ZѪ5��a[YL�q��	((�3Ee�Z�q��7v����R�_�YW�S��r�ƅap��>��ND��VX6_����$R�u)*�wH���k�)<�.��.�M�|�(�=�( J,���	w�Z0JG15���bӄ�z�BS��3�i M#~ϾmcQ�f���O6u�?D��sy��Va�ҖE�"����,k���_x���Ϊ� {dhx�iS%P�~��k�s�eN2�.yȉK�ļ��pńP�c��z�[ eĮjTv͋�����?B����^F2Ơ�ɣ{�>\9;�5�ىr�_L���,��}ӊvy(%�q�`�{���?9��+lzBA���[2hS�CMyv}��ݱ��V$#s`J�����YR� IV���:��8�7T�Ch_<�<���$�G{ܼ�5Q2�A3�26��B��ѥV�n��i���M��}b��_e ����0N
<�E�9�Ec�IBQ�F���|�2�/EP��C��\��f��75��ȗ��%?5˚�����]�z��qB�H+흷�u��s��0٤�^'���aKZ�qxE!�=�Xq�����"u�����p���X^4zT�	����&�Wk��1k�ɕ��d��Y�xA�3g�2]^�����%0+��/qv/\}���šHU�*r1LA�P5pN�0��M�K6S�`�����/^���!���D���O�~���)�E[��v���w�����ޯe�����}J<榰����smv�2E5��e�}�� s?$h~��j�|����6����>��>`�� n���Ts����m�lQ2�j�q��}�ۀ�<k3���D-b��l���#�d%^+w̻~�Nw����B�����k�d��Z����Nk��yФ�җ��І�o@0�ט���37�����7$�v��z��L�c��J�W>[d��^[p�%=���&TU�+$���l2�]l�\N���0`���aq'y԰����Y#�Y��u���� X�H��͙C=�0l�O�1;���� �m�Q/8�nj�S@�^�z���+ʳ�׆A �!��5�gZ�&�<HBL*��3�2���qTd<��ו �<0�H5����2�/�D�AؔS�Y o�{��}�	����|*�%��K���ӂJ�re,F*n������r쮆�3e���������T�w�!���[~�ͣ�Q� ��ԺCh�4Eq��3�G�JF��Yj5�pV��'�oC�iWV��g�ƶ'�\��$`��fո�'�؅�E@1ſt�Y���J����)�w��bs�4+5����Y$�/��'%b����F�f�F!�e}��\ <(�92�R_�&Q�4[��{��Fq��Ş�޽���M!�h�ܞ����"������1p ����P��'gK��5c�l�l��g�����.��l�;E��n[n�m����{�G O4�*��:��$l��`C\h�4;�Z-(�:*�[�PN��� �X^��wп�~��Z��`�~�-Eː8Rŷ�zS{�����s� �(��E3��~�L�i��R��7��>�p҃ ��h��=t�����/�@���4�
6RO�̔�uNo�-�\�xg�<*��q_��#7�z(&?в������o.�m�@S&��9Z�t�2hbZRh�+63����bɦa�����vX��]�A�K4��.<������W��P`��F�ua�kp��{�߱�����vl�9 �(7���c��,�*��]�nfJ����������	տҶ�4OZ���K��>�n� E}���wr�@\*�"��\P6�}݋Y^4�*�C�ay8������|�\[����)��[�����=/�yOK2ڃ����]��d�.��8?pOԏ�s�p&f�I��]����2O_��_?��a�$B|`|v���3mqO�%� Ƨ���R� �3�HѸ�0^���ߪg�b�iF6��W=�qE�kf�R·�6}��d�����^r��F���U^��>�a��q�rIf����bj���K�&�Q��H�*�����;rH�.�K��u��YO��V_RMXL�֒X��/I����h��M`#��"MN)}��+�x��Fi�L̓i�m�~Jm�r�O��n��Bk��
���]��k���?땆食���f���*<�td�r�=����+S`�uES����a��Ss⦉tղ���G����g,$Y��j"����!�j���	d�B�G�Y:2l]��єЧ��� @��=h�V
)s�2#Υ��F�4��nB��.go n�C�tD��[�tj&���ȧ�ܒfú��Nʘ����_���k�)U�Ar�Ud�J��#>��'\������)��'i��S,�9�|��t�u�q��.��%��:5��K����wGx_DF�%�_��<�&>��`73ِ���&��T��[�̇Ls�[zl�ՊK#���R�-�Q�KP��=�e[{�.�q���=�Ec�1 ��xA�m��V��v�� ��N�$�+���p��{�<M��oԭ�N��v`�|_�)��F��,��$��l�������c����u*1����9ܸp�Omb2�\���/٪Y ����y�x��[�$�(��E�8Ef���y½�:��=	��l �O<�̱-�-�]�D:�Aȧ{�\>�`�,�܈����r���t�k����Y��W��}d�|��4�9y��hC^��E�njU����e�!*�9�Ƶ�w[��ʋ�d@>�+X�[������sOB��ek�(b��|�e�U���(m4椉o���Zˆ5I�Fl�R��s���F>�"S�~,Y"^�A�o4HF���&��lW'd�`���;�`9|���T6�3ޥ�H�K:Lÿ��V��"�h>ƫ]x#/ \X������<�cŷy����"{�e&rA���ezY]����[e=r��;�u|��pz�K)��F	�U��(���_�7]�y�Oc���j���=:O��������B�)s�Yaܳ��5l�?�\_QwJwB"�y}7S�)/����S�9&1�Me���)<hg��d�p�mY���|dX'�n^{�q�Bp(�ʃn3sb6��+�6ꀶ�i|.��I�k�b��E5�Cb�㚃P�֚ʰ/N�a���8���*р���'��D���A���3��,����}���V|�=�=ﰖm��?�����[e9�uK�EFjD�Vx��}����{����FK��r>ɭ��GϠ�W$��S�q��ëXݷ��'}-��D*�*d�3kl�	�R��y�V։_a��We٦�߭K'o�i94�;��C��9�,� N�hy�]�"�(��Z-��찅x�o�%�D���T,���� �ͦ�]�UZ�h�ɿ��V�#���5b�Q������n�-���B1���'~�U ����#PZ\`a����G�5)G���U-?h��I�5�OL[�~��fUT]o]"y����|��X�ymx�o��g(P�~��g��Q|�<��W ߠT�dX��~�YC��*&�	�
G�^�����\-Y����g����ࣨ�Q�x�nj.�sD�0c�r��!�pF�'͖D]���e�PI8�躁���Za�
�N�ۓ��Ƙ'C����g��Vl➩1o)�� 7��SJ
.-AO,���X�@^��%��Zn�Q���N������!�S@��T��\�(��{ᵑ֬ȩ�WFA/�8ќCU=_�B�p��Y�x���Un�.��G�C�=�NC��}L�b������4�E�C�܂�sS*L�ط�I�������zz��V �Wx��E�0�a^!͝uO�3J(������^V���ͤ��U�>l"�T��FAZ�5����	�n#a�� �P�FNUQ�ʳxf#|�:<�,�-�J��wI 8�����PC�q:�������P���,=bM5�zi��_���le?OM�[���[�;M��XL�ί h���cg��}��C��ye�K�}�°W�m�`����6��$� =��e�hJC,�d�_�wF���pr�0�Q�8�.��]��RQ|��8k�/ EO/2��TQ/$���U��pI����ZR�7/�De���T(�^�e�#�WMg�[{�.�CBhs&۸p�|�_|�;����3�Y���b8��첫��i��\S�����)��Ľ�>ϲP��;Ak_� /j"I�gT89)�TF�?��5����%���s)���J.��b�_!���#��>'!�~�6s�џ��B����U�:79NC��W�Gu�����L�(`x�뎽if��=+�
J��(^�A���g
{O
��G�=J�$\��/^"�L!�%85ǿ�3��@��,���m�~�/�+����=�����q @��W�QPS�"c���֫
g˔H2kwiV�g��Ԝ�wV����Z����C�]������,��y��+dG�m���5nT0��)���r%mOkǝ��V�DwI[c�m{9Y�.�]��V/�����4�4���Ul������!�5l;�QR\1����$i���f�[T5}�Ԭɧ�tfF~��^�ؔ���;�,��{*6k�`����!�j�H����p�ܥ�d�׼@������l�v���'l7�mX:�;͊u�?"�R�6�3M����������k�Jͭ���-��d�����h�+���
�ql�8���%�f�EΛ^�褘�����U��C+pP\�sMB0���F��y�p�Q��	t�6&Z�,�צ�H@	0�0Xd����N�B��D�?������]˞8o��,� B��Dͮsu�EO`����G��C�������h�oZrj��0��Y�e����[���%I�ŵ�1k��n��~#aE�9��s���h�}~þ�{��-�2��P���<�D:�ek|V��}�c�A#a�)|�d=��A%c��w�=��b�]�s�W�1Ƕor�\�T�c�ۀ�@�VR�p��?Ð��֡	"�Ar̹QƖ�V��\��=�[��iIs#RVmx�p��E�y��ӎYμ%H��i靈�r�yD���߯B����4cEHA��NiR�}���䮀�� }����KS�Hs�ʰ�z���@�Ė��n�ڜ����up���ᱼ۟�4��p�d�A���^����� �Zi��.~�zb^1���Ŗs|݌��N+����¡+���g�ۏ�e�y���-cʨO`]����?^��X�N�3�Eat�fI3�&D_+�|">�.v`V���#�']���;~�4�M�� CCY4�
E���?���t�'@G6���$	��n^y)浭�Cw�����g'�7�h��ڶ�;Uz����j�x['OW�"*��r�6^�����>q�ȟ-l����*r�s�;�d��_kZp�ڟc�x���@��5��}�ᔍ&��������#�V�P��Dٸx�%Z(]}%eqH��9�7��$�v=��
����ݶ&�����t�P!��x&���,s�U蔐�/�3V��|�2_D
W~,��4c/@sg�h4�״㻈g�n��7Jӂ:��v}d��d!`-�[7�g�����[^�M&�2��D�qBʺi��� ������z��%s]Y�ި(<��V(�B��o�c6���w����@��x�� B��?2(t8����j�9��W�xC8G]4�~�p�/h��p�t��w �:G�G�㍿��[^�
6�1��m�XآU�*�/��x��l�L��p�Ygu��Q]��yF֝uP�z��ѳ,2 �E6�_Y��M������~T+���G�i0��|��@t,��.mͶI*���{H$�d��;���ӝ[����JP�tQ)�Fk�=�+пe�)#*aۯkˠ�u����8m�nyH�]�/|&�!1(;PLupy�K��\�Y�Pvx#mjn���)��}����B�XE�`^�(�7f�B7��	P�	V9��',L:W�a���ѵۡy��%~`��c����,�%Q~�a���~&>}�1򼻵n������g�Lj�Y�F%����.�g�'��r��`�
��E�3}����5��R�ld��\p8�����D�)ɴ�V���G|�8��Pƅ�0k���(ܜ�8!	�,q��S��k�� ~�K�`�ٔ��#q�r�ҕK4`�X����m:��(r�W�qb�s��' {,���EHu(����kR-�<�_p:��r��@����N�>G�cc��I"�6`��Bi��bc���'$�4*�ܫ�h5H���:d�������y욌�ȉ3e�k�C�r�=/�D] >�C5��֧�l�$ޟkN�T���dx7²�Rʫ)���9���F�P1D��2�+(�Λ