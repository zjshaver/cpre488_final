XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��2y~����	�\o����z6�<�_�/Eq��g�0n���T�y�}¨AֵLbo�%���7�����!�c�m���S�}�5����q�Am4�|�9���gN��� �輙�n���N,�O r���A�aVx|�G&����,�)�);�:�� -�10`��Ղ:�����Ϳ1�����V���ڀl����|H��ц��c�s�S��8�#?��m,�����9��vi3�H��?;�2��9��\'���J&G�u�)Ih�����|��u�c� :���;���6��'߬d���d���#c����\^�N`aJ�.C��(~�yp\�WR�mV�ϘvnJ]�f=-��u��l�����֠�C��(�����Z@{BkM>�|^��i'�l��ŧ�^��?M*��l	��i�%����ω��Ch^���a�7�mV'�0�k��^?�Ҵx������Y��QZ�G}[�B�װ�h��]E_)�eS�� �>����y��D�����U1�:�Kg�nFZxX�[
>�k�Y�-i8�s.��{��w��{� A�����"*�ņs�)'��O�$���5�/��a�͇O%�)L� s~�%:�+��x�%�y����K�	,�&�I���˟K[��˥ơ0S��u����p�{�.�-�@���L��v��L���W�$��4Ѷ2�)�r�9$�/��V���։ӭ���䳗W�<&&�i��J�>vb�Z�C[XlxVHYEB     f9d     6c0ۣ2&A���+n��v��z�4�[��x��r�?5(���{�b��L�\�RM��	"U��מ�У�A\�_f{w���]=�K(���C[�Z��A7-.è����fi�����3mB\�X� �o}g�vl�;#������tn2
9l�Ir�ʓ��S�̩�o�Q�)Y����-��m��U	Lf�If/3��L���FYt�o��F4P��wy��m4���[�wr�f:QiAC��1��0�3o>=���h]9&�ݡ�c�K����߈�P�A��-]/��ùѢ�&D[��o!Ň���g�:�Yo骃p�"UH[��
�s��ы<������jHǍ�?��?u�'��Qt�"�w���䍉&��X����49h	J�J"�^&���_9��=˺��=s�:Sa3j�#���f�����,��G�zKb�($�����@=�u
)��U=X=�4�Ʒ�: �4羱*����ޛcgX�~f��T��Tn�����Y�b5�h��N�#�B�ޞ�Tt��D]P80<��w�����Hʇ�CF��'ay�&Ph8���)��߄5��YNFm5K�rR��yN��Ӽr�����|�|��d���5(ip�/�K����)����M��>���r����q���Fm��eș��5͋Ez?ݹ�D��;>�X܀\�dt�qoB������B���a����8�5 ���Ԣ��Ig�-�C�����^�r*��v�"<ߏ��RE[ǡH��^p�,X\�U'?�-"�=3
6��`9쫤�md�A��/�x�O�H�ݧ�X�Z:(�هb���7�c��G�Fw�/�\F�P����SV�v�;���vZ��~��c*��j#�Z!b������2U��������D�$� �j)X�ÏՒg�3^�� �Ws��e��_�M?�Fb~Ȩe��cDC�N��F �
�)�L������18
m��a`��]n
��?
EW?�U0��컃ˆ�֠c��������h@!7�l�P������ ����(��^װׇ"��h�
�I��`�������5�iq�R��)��K��7r.���~��; ��jrM�3�_�:�;�MJ�w�<4������ř�oM���0�����D{z�4)H��6U�'�[v|V	p+�7�!�f=ػcl@7@,u�P�O��>�|�����PSK�x�eڂ&��3Ч��Y����89����8нr�2>�iO�Iz��-x�-��AlZ�[G­�^�q2vφ���`Ʃ�"�6Ji������pH,�vMY�P�7�v��YNwUL�j	�FGy���"7$�g���Zh�d�@�	�+���V|G"����J�%;��ۋ�(��-�����7딨�݆�8� �#C�Po���@����4�����_Z��;��F����$���J���X�i�J$�ơ�@a1�Dג��$AZ�2v�[asBB	FM�u��u+�yW<�6�=❽(�>�����h>C��{��_zq���af�=;M@n=h/gj�𕶨��-"��d׎�O=E��ᰲ��zM�#S�4���';�{aUP��q����M��X��x�W��k�h�d�+���2q�ת��C�DO�6�	�=�Z=M����E���8^��jx[�n%ul�S/�I���>�25��U' P�;��� h�s�̥Z��̔b�S�%���_�-Y��K�M���u