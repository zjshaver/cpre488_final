XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������N�F���rzt�z��2���������6�?,�b��)z*��4���VwdA�:���;c�TͤD���[gP�m;xW���a��X�� .�nP'<w�_��N>��&��+�f�~Z��#'�����5���!gD�@W��{�-E^kUe���Qȡ��8�a&k���~���&&F������7�E cȺ�NU�s�M����?��n����'��������od�0X�hB>��g���O]�Z�\F"����0c����(o�=�{��t�vc�O4�q|4_�ɐ��:�>g�����odi��:T�ՄR���<�^��5Lc�{!8T��O輳-NL0��͐��i� U��%	@2�7o�DL4��s y��h�2����e��H�p^�gB�R�C��;��5�\S(JQL�������V��)p�P��'��!�&��{!0�`-[�*�9%T GME]-}�2��&W�nn�����"*���1��x[ӿ�&��G�p����d�sL�k���L]s�M�.Ңw������Wj(���E w��>>�{`�I"��5��ݸ/s��|�������9�O	�]�B9`X�A#�8L~�:~gt�NL�;z�7D�|.�~ڑh
�1~�L���7Z�	,�a_����H�֎�ALZ�E�G끴J���X��7���Wr猙�!��J3�?��o�g�2;��Q���]�}	��4� �A*]���4���ꫪ��b��XlxVHYEB    fa00    2040���a���?�������X�.!Zw-��*��U�wd��|�,>��,�׳�yI���h�ܼ�+�t
Z�����%fA���Ix2i�L41�%�2��蝜�����MK��7�8���OO���#�o��ݾ���V�[�J�f&G�Z�`�=[��=�ퟨf[�M�v~.�}i��L�m��n�w�"��_ :�7Y���@��ڧ1>'�����-�7H��.�k��u�k鼴F����nXYN�R�3��Si&��x��Dn��]���v-یX�D�������D��Nu9?��Fz�YN���x�():�o�`�#��yw\S�@�L��W�I����qL���J��"b�Q*Ͽ���0��a�RQ)��C&~���x���͠P����-)Q�.ΓT��Lu�2H���M�3�
F!/{�g�b�Cԫ�DL�Nh�'���� -�y�J�Q]k
9��3t�_92|�WmY�݉��g�L[n}'�����B#��	�~�iLN�9��mzGU���b��Y#���d��2'�p��t.rm`���w'9��<�o��T��Q)V�\{G���_���}�Vl�\k6��#4x���uǵ�B%.��<|XTKJY���ɚ4���Q�(��p7���8[Y�ɤK��{��,��>�C&ì�ٯ��t���h[����n1��Ϭ���#���B������Y�<�O��[n�}�+�_�繎bp����҆�ZѻVO��aʜ�X�E޸[+�g�X,#�[LvN2h	�����,���NN���0�+���OJ:CQ������.�|�]D��g�}��>}�����?-�>��L�{���РCN���؂Ь%��|� 18v%9LU���0C.ܓ���8NB�f�l5'����@�^��j��}��>#�&7k��'���\��oK1��z�&�)��bXܪ��R����l�*�� �0�g�Z�m���}p�+*@��=8��L*����(O.�E=�O���������[��"��/cpϑ�s�J��y��1���:L@몶7�S8ʫ�I�Z���J��ׅ�Ѱ�t&dNOp�gK��k粉��u$���t����S�G����6�^�Y����p8��/EJq_�@�Q���Z[G6�4p��A�s���uH-:�*�0�<�_S9����7UO
3|^݃4g���ۯ�{�a�Lqwՙ���e+u6�O�Q�g�f#�\)�/�����t��eO����]@y�l2<Ӳ|`��\��Ӳ o/-�#O���9�v��Yt������Yp�xWch� a��p.�3a�����4�pF�~��Q��zOA隔����X���hh�匳~�A���5��:3F���V��"ݫ1Ԙ��X����H�P>�ڱ1D�`��,�����8������U��~`�I�(�q�*��cl.��pT��r�9�@���DDL�~E�����$iV�w�p��Ө�hܵ"�I�9_��?i���d�J�rMϲ�W�]��.𸝱"�� ��iy�O�:�@`Cc���!�ԕ6�	��z�<��R���ePezo��nZ�q�f�qM�A�����=�|�L��	T'n�㚕g>��F�F��*�Ƀd�k8^���l��ź$j?���A�c�Ӆ+:E���5t�ZQ?���"���h���GA��5�)J��'dZN�:b��	�e��H����#+z;)��=�p�\���G��ݨ�vY쪁fI���t�z���5&2�� s��|�:�1v���e���R��я�WV��='%��:���>z�
x�m`�� �E��~C�ٓͥ`=D�;x]1��O8-Щ+�݄2��x�QK���7��l�	�'w���Ӫ~w0q��`g�*�h8�c�-{�Vm�~WI,<)Rco1��U	�Z&����hr�9���>3}oødm�F$ON�o�+�<c���P��^��ڃM�U.�ߗ&ς�<C��k�;T#G9������YF:�1:�����@w�e7�Yв�ҎQ[8 �7^G�S�ֲZ�JxѼؗ�c�����wX��f��{^�v�`���X�E����p���댉��Dtn�(�����zZuɉ�ޏy���?�`޴��ԩ.0�w����t5���I�3B�s���"��x�-��}�ݕ�,j�s����k���耿
��/ܶ_�T,���[��K�����-���	&=\���57�Y����{� �.~����I�������.���h���H��/��G��pY��lW�GE�9JzD��Bu��c�_�}q�8ռ���6�W�z�1/u�^�hU�����u/�OV}0N��h �j�?ZӚ�-|5�ǹ���o9����B����o}:� Tg�`W̨��6Fﲙj�mMr]I���Z�}i�q�d�r�}���X��V���v|=V���I��?������ݻ�4��VQk�l}d~sL���v\y�9^7{��̤!h�1�b邜A~��0�곑����[���D�Z5ZRG�ϲ�gc0� �.�Ro9�m�~�)�2�깉+s�W�(%�yH+���[ǻ�u0/�C7���\���R�}Xb�E9�]�@3�ع�r��C�/��s�`�:� ��M��N\��>u =}��]�-T���8ɾިVm��Q���p*�{H�!�� 1������4S����t#�7��")��2���\��� �	���o/�_뇸upֱ�S�){�c�5�L钝�a@6��;w��)���@���%-�a�Q� ?m�jMn�2����=����[qXjˬ$`T��/A�L��C�r%�M�c��_�CXr~��G���y�A^}G�R+p�~��}Y�|�h��U3 >�A�bY���$����0@
�E]Qca��A�V;B�����:���}��
7V�*G��B�0�]�.�j�?��%%���&�is�\=4��[�H'p��z`\�7�@�ݐ-J�
E����Q�d����[
��t��B��m(=��np�����T��~kA��%�F˜��"��㠎a_2�a�j����5��Zޖ#�n籺� 2<(u�x�O���  8�?�'s��K��[���Aֺp�ks�7�及W]�$A�	']kf�������.���X"r@�i`K�ʴS>[���V.�!T4�p����fxv"�&���rd�x̲y|q��v��Ti��S�<�%���/�I(*���BM���9�p���	����>�*��Ô�,�UoF�,\�aS�ws@��Q�9�l���;�q��l�)�.��>��=���?�%Z�N�0O��9��N��S.�ն��ǣ/cu��p�d����IZ�Ԃ[��>^�h�!cy-��6
e������{8�<���%��ǈ��5�=�,V<�T�_5���+�;��^�����C�sqxќ�&�>�<R		��Q��}^�k>���]�V��Z�[-T����k�y+n��r�Fw�R� g�,�]��.�S��:�!җ؝�b.qHЭ��om��Vލ���|+"tL�뱬AI@�d��������7����|�m\&j���R���`�?�>.��U�vu}�һ����k��#f�L��?�`¶2�Q�>*9�b&gñ��H�����gS�QU��$R��+D1��B9<�E'	�f7���V1C��(��f�1�
O�	e��3�E�;6�ն� v�^PrSAT��Ca���B��a��"�$=*����{֕�3�ͫ 6��hȆZ�����R�$e�{���dpFck�
���?�����Omd]o�h��	���5�
�����0ή�ˇ�t����Fi�ޝ��d23?�C�N�&�vC���)l	���,i ��a�������ڊkCj�8Ƙ�ē=���P��ޞ�U�GL�Y��Cӊ	�f9ȕb�
�^�(��'�2?���I�U����\D��HSV�k@��&�����p�	�PȔT��t��ϑ�sf����"�N��2C�MFI�-0�O�=�B"�)X8�����
C�<�G*=��#{�Ns�9X�R5w&TN��:Ed��u��}-�fB�^�d���K��.���qm���q>%C���N��!��]�S����K]k��	MOk6��z��ɒ6�|���攃�̋�*�t ��T�
�<�م
c�*d�U8�ա@�=Gm������׽��AX�a����25��Ai�or<�p\��<�s�4�:yo�.H������OĚz�Y�#7�΋���{���
8iN&8~m�"�4�YV���|J�C��,������,A74�倷4a;T�ǐ_����\��ӵ�Y	qVt�B+7��B��Z��o;�O��� ��IU������j3�r�~����C�S�&���ؕ�:]q}d���)�t�_� *u�����%�rz��@����
x�K(����B�Qڋp��L�$�Fyt�l�NPW�C���x��<�a90Z�3�ThV�+[x?6����ٸ������?���&����?����^ʲm����M������Y�d�P"� 9�@��},򨮉6'V�|P�RFc*#{^�:Nڼ`��r����QYf�1�W�vJn�ʸ��/�
U�X�� 3t��dgx���ŋg8����Y�O^�3ߢ�Et9}�s]Sr=z&,AL��|���Z0E�l���#��ƿ$����xU�^3�]s�|���=���~��oxT���?��H�wn�t���	�͍C�0��Ƃ0���zn�.+��TB��R�G2�k+���41:����j����4����M3��}e�xo��>k����x��D|U3�k��,��q�l9�9��JϦ��|�a�/,�8��0^���s1�3	����#v�ft��nS=��$�a:b/�L ���U�BĨ�����؈��[�uq��*��M2���z)K�Hm'�p��XÝ�ۍ}��F�f�������CхĪ��#I��h��ͽu0R��_��>ۿ#��,Xw�ʂQ��<���H-X�K��@V�zP�;F��6��e���a엒k�2�^��s�b��?+k���,j��U����v#@�+����k35�Y���W�m�=�0x����E�(�q����H��㜩*x���������2d��:< {?<)Y7<����j��Jc�DE���-��<ǿT��g���[Mל�pn���������/L6&^��>DQ#�\9]F_q3"�T%�^��?���C�ؐ���3���|��.NB1�j�6�3+�
�ى�c����(��H\�s��[��]�o�|Ѕa��o@oρcwTb^�o�A͖m%��n�%1�Z��1��\߯sgm��R��P�{�ԋ��v��/�OE��0��7B�8��}�O(�z����S���o��I�%�͢1�Z��F_,�_�x2��w��ׇ&D\Qَ��55��\�A�L���kIy@�$�^x�S�dPY���w�Na��!Q�W��(
��$՘�}���C�FE��^�bצG�����:��|�S�Í�r�O
�K4Jm��r�r8G�Q+KZ��!�KlI��� ��wXYG�x��zZ%��D7ac������Y���|Ձ�}�F �M����A��&�{���J:H�ܯ�?\���rԤ�U[��4�f��~�s��g��)+��n.�h������N�#�:�l�W���M�^��Ӆ�����),�FZ<��j])_k���F��Mɍ(u�Ѣ�r�F�u�ٱ2L`U�?m�'Q$�p7Y�ƽ%~,��K�>ε���E@��Ѯ�[��^�������c	��k���f ��Mv'Ɗ{���$j;��g�S�y���5��$\��T~�p��w���Ƈ1�@��y�)c�k�?����R������N�fK���r�491�U~fr�v�	�Vz�a�p��>���	7��]rH�6���HV�z���t��r�ZN〉����g��=m�����{��L�&�+�*:k0����̲���=��t�x��pE��6���e��� �;dl���3Nq�p��:��Op��)X͉�4q�zfT�'��VŸ�@�Ҝ~{�X̒C:b涼�����$>���(�5�ט�	�h �{+²����bx���`"�o�Rgf?݀l{�=�.�[�d���Ɩ��\Re��l����1�0��U����ȍ��ws�lu�<�+
� �.0��IN$����D�RWB>C��6q?[��v����z��M?��.L|Q��%}2�O���U�怅�d�<e4��6��9x�v�:F�*B�&G)z�#�;^��e�ҡJ�*��JF��f� ��K��ůmiB�>2@6\z�Ql*e��]�[V��� q��@������)�dC�� d���a�m�Pz��7 {p���r�L���-&���������|�^��`�mjA��V�k��n��h�11�.�aCH�P&?�nT�&�0��v(��
v<����X��Pu��;]ѡ�׸��fYPC��2�%.��0L���R!�M��(�o��ֿ-�����Pg��	�����j,z7)�4���bMu?f��C�H�Qm�!�l��p��CP��qJlx��o�F�Ea�yE�.x.M떈��:
��֙��	C���u�����*Я���e*�3-h(�F��޾�b2����~��+�#�7͸����Ե�(��Uj+Po��@'���h���i&��9F-�7��_#7�����U����SeU�,�8PT��SM "�����<)�ς�ϊ`�����g�$���^r�%W�6����b�ȅ/,�N��Pe^ŔR^38�zOp��Տ��/^8�n���i�4iT-Z�h�q/�G�6TX��Zm;�_�[~[٪ _)N��Æ��1�߼ɚM��<?,���菾^@uoth.J��Uz�&"𠓫�7��B%����8�-��4,���nt5�.�R5�ċ�'��ɾk��m�af���F<Ŭ�(�����6��<q�Yww���t���YJJ���7�~k�N\
q�7tu�^BW�}�eX[�oG�Ԍ�j�PvwF��?k&n6W��:�TN�[���R���&��-g��#��
���g�YC����SOS�o��
	Qߨ�������^f�X�Ǝ:uPF��;�ܤ�^*���ȎV!L$�EꁖQ+N�пS��`"���v�ⶉ.��ۣ���:����˓?�|�w����8bZ|��9��W�Y�%=��z ׁHvg��=���]�s�c�s��N���5:=��F��W�y���=���X�y���Ra�]��xDŐ[��=V���u���zV�wXd�4�2"�O;/7
�r۝Km�9�ּ*��$��#l�S�����WER��ݪ5��i�4k��?�\gU��]�oE��j���ni��چ�'}�M���d͞��&�h<e��1W.����}����-�Nt˥��+�[!
?Y��S�7��3����=t�C'�u�q�h�C�EH{W鋹��I��k.��ղ9	3Mʜ�"�񖾉o��d�4�/V�م,#���D`z}9�b��B�Z	��Մ���W�x��w�|%ܠ��F��R��������Z`�cyH�#�v4'�g�d��dǣ�Z(Hf\�/w�P���h�����>������-�t�����9�P2h^4/�/�~w�v��݂�S'�̀Ks�v�&^��L�����IYX�=�c/�p���Z�G:��s�[��ם
�߷cAU��&��p�c��a�Z�J�ס���)�b̻��/���2��M�w4U���*ĝ��=¬���RO"X��!��rߋ�x���z�)�����5K@�t�*��HLu����a_��l���e�&��<?z�I���U4O"��&,LHy��^)����#s]b��o*"��I��Á>��ѓS
�4@��1%k���MxϬ�K�C�qOF&�m��*�bJ���j��M����fNC�q@rjų_�m"e�*s�!0�I�7qo�N���*�?�L&�(ךP�"��W�j=�+*h����vy�qV/�ww��ٵ�g��7���y���S&�#��{���]s��d �5 ���ֺ�&C�L)���2C"�j7'��
--1oXlxVHYEB    4f62     b50x>DǕ��[BP� )�qv�ra=��X&�#�94.�cwN��f�����GQ�}��	���ߧG�UK�r�p��m�>'��a7W0]܅�:0`�ʽ���'�w�V[�Y�+eQ92[�ӈG����^���(/�2�s0s/�a�{���T��8�|�k*9�!���4˽��r�$l,��P�U�"��B�o�1.�rń�1L�$��Ԑ��/ϋV�gh*%�Z���7�A]��@������{`���W�*��"�mNԕ��-�@��Oj��w���:횶!�sUs��-�r0�hI���1�Mo���&/�
172�f#Cb�x��C��ۍ�nd�!���z�c�þ#��&��3���!�������*6p	�:��؂3S�c����h���H&�4r3��Y�A	�sj��l(}�X��(J��Za���p�� �8C*��v�<9��>�m�l�5d|`B��y�e��IQ�R��Qm8��ʘ����H�����\�D�����T�K��ˍO��&���S ���	��,���ϥ�I���+�D�����h	�an0��ˡ�8~屝��L�H�%~�-������?�˝��kgH���͇~��g�W���u&{[i���(��þn����UQ��y��\�冻VՉa��#X.��<��+RZ�$i��:ow�꽭�Is��V����@�[��Kn/��$Z"�!�ú�M�`Sx��g�(B�����`!��$��2�9��]�0�.��a�Z�ܺ�Pz�ۗ��Uu�} "iX�,�/��~O���u�cu�:�b;h�!4�R�V�+�P��&^��y��F�l3�R�`o��	���#����L[�NM/D��,��Oi�M�"�_�ߣc�-�a��n��St�p��y�����2H��%��}��LR����Q���u���Z�I���4���q	/�L�̌�C!��ϻ��9�k-�,���<��,e�9>�lw.{�Z�����g����fY��5��$������d:MA`�'ܴmv�
���)��gZ�cp����l|+..����I�Օ�����ܸ���@�P��m����s5�)��9.�N�f�La4��*��ȞT��X�1�H�[S.v|��R��C���<^J����Y�����<!����)��"Th���i*	����a�n���(��C�
�۪l'z�Rv��:JF#�ɩ�*��/b��xq�^+{���U*�0��b�cH͘_A3{G�+G���n�s�"�t�G7���O�Yk��������yBW���w�	�9�+����-���!�|B���Ⱦ��A�ݵ_�v�N��@r�씽�1����|�#k�T��!tj2�/9�2M���wx:����6&��a�l&��G������?^#=x
��p�VL13?��Z9��w���˕���޺��m�RRn#���iٱ�3͝�Epm��JN{aF(G��£c�q��j^jX�����z�Ƭ,��7�p�6�Y���M���}\���%���}��Ⱥ>r�}X�=O�b�Cs���T�	)9��������e|B5��)��mP����<�:i���1�U���*��es؃VZ�X˕�sK������n�m&�#�;�����B��kӼF_[í�C���kÕiZ���VM^�����Wѝ�>�9W���v��X�"#��H�����s�*)���c�Pk�(�Mz�Ƌ�1���x`��;�:�F *��(�),�F�w:u���1,;Ǧ���A��Ѷ���g�WMk ꤶm���8J��\]��1C;�@�v�aZ+JF�1�溲b����0?KA�
6¡ɦ��C�`�y+��|]������Ta���m��v����5�X1c<�]��	;�y�8�[9���V;�X��%~cdn+Aa����)\	�Z����ϊ-��ޙ[gܷ��_(c!���ZS)r�DU@~h����na9��(6)s�5��,D�S㥂e[�=�F�N�byS�c��1-HT���z��Y5t,{���7Y���Pc�cN��ے2���@���[��ŀ//t�95�O�[oh��0�H����R����v��GI�����z��2)4E���u�������=T&/W;�^�~�!��;&�������1���u���a�`��𺡾y6�2�=�pO�lT=�,�K�>.`<�F3�;w'"�lP�K�����E�8�GVH���!*�s��\��	�x�F�W7!�v�Vq v#l\)�M	{>ź���L��D���F�T��b9���Kݺ�|��z��5�������8�\�|����1f�&�J� B	Ǐ[Z܅��<1)��ȓ��i��#xe��� ȮP<���u�pu��	,E �ڍl�����I=_/tY@12�|?\9�7o�J�� �֨N'�^>�{�gte9�������lhs���,ھ���3������J�3Ǔ��܄9<��x�Y͈X�%NMLQ�o-���K��6 �s�3�	22j��0z�V9*>`*}�P�:�R|	��ݦA����	�p��}pq�`��V��ܘ��rhy��9O���L��x�u�����ѼT}h�aF�sQd��3��|H�v@-�+_�/(T|z���W��2�풝�y�MV�7�al]6����]������1�Ug,��/vO�̯nIˆ����[ي*lX.�6.NYb��&����&w�X�2&�+Q���Y���5�ͱ��@ZO����^{���U:�+�k����f��"�� y��w�S�hF�"��pQ�	+�4�_箷#V�=#H"p�3��E!4o�	�����z����K�\)/��!u��s)sO�mԸ�Y��