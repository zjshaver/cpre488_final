XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������J�QlK=I�;�����~������ה��n5�� N��O\��p�U�m��Syo�	b��S�Z��=�.�j���{6J*{�ny{��&q\�+��������u*��w$=ˬ�k�ꐒ�����ޠa�G��TW��Cb*��Q����,bA���>D�vdC %�~��BmU��'*P���>�d�E�(-H\�RG(3��J{e ,z�^zsPW��}�x,���Y�W�:$�R(�<�'��\اΣ ��1>$_4���Ҿ4)��'�H�(ܑ�Z�00_޳�Amx��8�9B��E^Ff��{�(9����n�������20g�}��j�0�rӖc!�b���כ�	.�H��l�{�2c-�q7�(�.��b���Wd֊r�#}�m>����۬`9�m��Z} �+�(qk�d�'�\2-O-���������fA���*쓪[*�	.O��R�s�_�:��U�m�uc�Z�ס��OW��v���>A�Z׵�5���� ���@��3Oց]��E�`)��и�2n>���\�n������S��C�A��@��> (g�2	@�5�%d*��"�<꒶�����Ά���s�\�N���A[s/�,`D�#�����c��Qɮ�_�e�#3�Db=9��i?wۖOt@y��XC�=hY�Y���Q���_~�d�֥��<�rUp�A��h��Ja�󐝽Ǥ���pZ����8-��&�O~`<������T)�*�~�������9o���"���*�f�17ZXlxVHYEB    2326     980ԕ�6�]�8B:�b
��&��P/���R��-���2[�����!�ϣ�CY���,��:���*vb#d��z\`!���6w���:y�����K������Q�I�����Θu�+Ut��Ɠ�[j>���E�$�w����$�.2�Y�kZ�Y���@f�G��b{-�:�M ��|_�)z����tF���b@�Zbo���Vx�W8���ΤEm�b��_���j��UAx��O@���4����L���O#,MZ�p�DO�FIZJ����]��=� ������|����GQ/Ҍ �&t?=c�����0ݎ�,i��[�OM��� ��W<W9����67����옗���/V��;1XQS��ܜ�o� ̷	DѶ�{H���VP]?��#EWP ;�I�a7�z_�P�pۿgs;��T��t4?��E��Xz}�GcC�K���� ��n��$bUſ��Z�^�_���d��2����'�.?��尸�( ��Rx8�B���oyН��;��f�%���s���S�T�1���r�h6\�~���f��a �����a&���m|�̕��ϋ �};�+�^���(loY=hQQ+�n�O�j�uE�V��6���{�x�O֦� \�an&1�,��pʮ���D��*���/��n��u%�A��g�T���	87Zo�t��#Fn,����\F��̗���W���;u֩��[���˅�&9�??l��k@#�C3dta�֞�(qHnt�t��Da��(g�c��9�"�q�@��ȸ��� ���j��s��\��{��vQ?Ub���/�cdm�/�L�*;�$ׄ����U����D����
M�ѥJzH&�dH�)���k����3�PH��I�\�B G�W=�?}��Ԃ�E��~�}Ij���&-F�.=����i^�=	Z�ڝ����\(�}�s@.%&��޲�'v���ʼOA�ȶ��=d��Kw�M�1 �-�x(��P��G��#Y䷤��0�y�eV8+��c������垿l�	���������#�bbB�#]6���RXO�Gk hP/�������su�(�Z/���;��aY���_#�5��蜒i÷���<���K�����w�^�xT���X�8G��z�>	�	$�!`�yy��� �EԦ��^
M �G���I���j)��ԟ�b�	zGkD|ք�G�~-��qm��'�Q��g���EN+y'�2g�Ƨ&��v'鮼4�a� �مxi��<'H�3��Sm�
%�=�1R_n��@O�b*_<	]Z�+�)���K�y�!�T�7�|�p�?;�� ��FaXk��+��P���▫NH�6��>�}�U4dD
M7yG�h��X`[�]B���F�	+Q����m�U!�I�`����A#"h��ټ]}F�P�w���׋5�4	���çp�Ź�!	_��l���Z��#��*�G��gZ�B��E�P�J�K�&��`�̀z�	�ƄqLvR>8�2ȝ�7�^{�������/�k� ��A�Ƈ�;B*oidd`؇,�9�+hK��o�V�6�=�;9ǻ�a���\*Wv��{�]�U�<{�fAlZ̶g�.��2��#@�~�\��X�<7Z��*��k�&�M��M�f��R,:{3N�]�P�~�   ��b�n7����!�r���S۰!�y��X��ܽF�ދբW�2�i����a����*�W��9�<�R?` �
3��A��os*�]p`I�ˉJK�v	���G�Q������f�����>���j�������(��I#>;���]&�����"�����6�% 32�{���ϣOb�7ع��]Z���L�����a���}X�f�3F���Uh%�x���14Ngw��Ğ�=l-�Ȯ-���+�V�}�����?*���@E����:m���ϢL4�-�� ��}�R_�h��F�ģ�J�!�PV*�s�Hn���,xU����Sħ</`�l'�rBh4=�l+�O6�\{l-��3��9%��9�Me11��M�T�����Z'jE�kN�#I�@">Xc�ŵ��+ytdә�!�u ����{*��\����Ab3DU@ɨ�~]"_�\Zχ�T���)�9oe�*�S�W~$h6,:��C%GF�"Y5�v^$��^�D��� u
�X�,�(qC���o�6�kC:������<(�/8>���7���'�b�8�����Q���d�6�3�h�h��4��Z?�]��rV�Tͪ��ӳ�h	�������rZ��h�[�����~�1q�������΋�e�yjӀ��7��@�����i+v*�5���HL�N�ĕn$� '6U"��ĀC�j�1N�h�2��R\�b��>�D��ܯPIb�>�m��v(b��