XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������2�]N�0�=�ͫ5�v@�kG>ƛڦ��	�Yi��R���e	iM�5�M�TSO����wIG���$סy��ߟ��5Y*�����y��k�3K8k;������3�C�r�~���&���F�~�N�T%r)�+�K���8�6hU����Цgt�;����1df�g,�Vгϸsy��.S��K`� ă����Q�}'ㅱ³�\옽���u1S2~�H�/.x��j�i���Dۏ:u���~��ٶ��H���x�_�w��m	�A�?�����n�j��'�(Щ�X��������L��8r]R,lDa��z����x������*[W��8��o��i�g��I�}wm�S~�8h�њ�`Q݋�Єu�^��* E��H��
�&-���8rV�Ho�>��p@�o�o)�;�Վ�J5���	uO�} 'ed�@Z������	n��;�H¢��CoyP�K��r��������G͠	ϣ���Ofq��>����F%S���C��$��-L���F�KS�*8�|K�k�[\��G���z��*Tz�ټ~��{�(P�P|Yc{���O�HZ�=M(w�bP{oAq�6�,�����dd��Ԙ�Y��_s>���ڎ��3���/�Ӆ�ҽ	�hiz�������O�Z��LS��E5)qH�Z=�?�+Z0�����rWi-S�h1g�MH�@R� �KЕ�%�� D�J���Ҟw�v���i_�"�EUn��x���%�-
�+ˊa�XlxVHYEB    fa00    26e0��m�G�1I�
�=����h$����ґIzS^�|9�]����w�&���mFA�W����(�pC������Z@u��"觴�����;�<�s��%���:.w���:~�J^�Ƭ�l�a9���0�TB�$ʩ��Ѭ)e�|Β9P�zY�̮��Q���f}"�K�2��p5��l���eч��\��G
�Y��J�(����,W8JB���.�A�xބ�e����.���{�w)��JRçA�m���!@p֗��c�z����{9��%��c!l�g\.__� ,�]#?��I��:6vV��&BC̹�Ʊ�Ns�%���XX��
�������p������{���~��-�%�s�'��J���p� |rc�An� )�M]�Fb�-���a�y�����;h��Է�Nlᝠq:��K"�V�wz�%�E�7
�����A4�"5�G��j�]��zN�s���7
3A�x" x�&R �J��K�X�L�|�u�4��*Td�nC�킺uj�L�9V���(%�y��#r���
�_��E�M�IO�f�����)/~�f�)
�����i� s��]l�������,ѮX��	 �2�x�f R!�O���T��JA7,v�)#{�����ڻ����_Ajѷ��}Gt�i�s��_�'#T$��1��+2C�M�$O<����2��_�+��ZE��V#�aB�<7���.Z�i���5�Uku��J|���Q�3�&o[�߀B��U&A��W����h� �}Ӌ��KW�[�i��&������[�`2O�,�f��"
���&�����iV���.�a��a��l�}i2d�J��W';�fK
ڠ$G�=N"o��i11(��E��^�xܨ���f��*jҷ�VN|�E�(��w�ĚB>ŭ.* �h`ӡ�VY5���a��k���K�H�^�-ݏ]���$Ő�O��{�t���cVc�_�������D��e�M��/�hc�1=8����I�գ�ĉ&��p�w�j���FeO���GpЌZ�&<�/ -H�<A�?����Yb��UK�v��Hk[=$����r��7\ވAg��B%�3��K =H0c:�y�Ƞ�IC�k"b@8kK�A��v�&8�M딭Vj����a`��X�-��IW[m@�Vg�\hB��F��n�lUOr�?;��\P��s���/o�\�Oo�=>����Ye4 ��(C#�?ئ,{��fI;�������A��H�:�Zr���ŏAH���m��[ �9:ċbD��L�n����>���-I-WzR�o�n��NFC�df��8J5���$Ʌ��ؑ�G��PW7�X@s٫��/s���W���=��1hj���z��Q<���.G�O\�Hf�L�xQ��/���[`5���b<ہ@m(��?.qs;����'�I�
/V��ǆ�*��+���0`	}{x�n���f��%����"r�Z���=~r�KfB}]vp����\�ڽ��a�a�t�>��\f1�e���`�#[c����M�f���װ�%j�Rg�C�T-0HC(�`�g��w���J�>y��Yǌ���F|F��fK�h�[T��:�ˎ�Z"V�ǃE�B��0�4j���E�t�q�����1��5��dO��#ek�[��l}K�bI��Ʌ�#}�䫮����u�p�#�C�X2Ǫ�%A$v#�����ė�qݱ}��T֏?~����f��@�a�@�]�sn�L`kς�C�,\�Z��b�S�R���tXG@|W�T7W0���*�)Y԰�Q�F�c����P��L�1%>\��a���`�|o�\�5kz�zr�I���}�E�ᘠ݉bl�F��&���1�4��� mw�@4ű�H��ݶ�~cy��![���Y�� Y�G�2j���^q�V��ؾ�͈-'�.C��I.�R�:U��G� �E����Q��)h�T�Xteѿm?_��4D���n����ta�GOB# r���Lq��QʧO��Za
y(+FP@ ��fx�"�'��'0�A�ɫ��$i�>�j��?}yJ�W�A���Q�v�FZ"�$�^��%�
�_�����q��U�Q�ٻ��n�re[�C��/��L�{HI��6+k�~��K�C��uܭ��qA���7Fn�:�\�,D@c PS��Yd�S�w�?��?x���%ѭ5ք�y%o��Q�+n�.�}��3�0X��/�K�y�T�.C���w��RV��������I���ͯ�^�əYe��Q�����}7��tϘ�-\���]y�i:��uƎ����WkY��q&[�y��r ��I���������r܂���D�␗�pf�����m"VOj"�yP��\�r���˳M�j�|�*~`jAk�Zr�t?��V��6X/a�S��o��*�=�=�ތp���7'㙩��-��<����^����t�G �#�Ҷ沘��*�F�X�O���O�M6�Y_��'���Z��T��+�o�lU=0@||k��"K_p�i�r�'"�w�"R��Z��>�%��yϚn,�rI�h�r:�a��=j�T��<~��c�:�����7l���'��>��}jB�y��MQ��9	b�ћvǃ�3�
�r~%Ÿ2۬��ҡ)��h���n� �z�gH�������hMuLv�ME�(9��w��QU�g���)-���z&:=��ٵ+��瘲d��';��$^g�����
�;��U�Ҕ²��H�5�ꬩ)�63�y��}��,�w�z���?%���+63�t�7�^q�i�"ۆ�v�S�F4��3I���v���,��(�1J�?~����b�>�|��P6��E/(F�u�����)t�7I��H�B�'�;L�YJ@�(t�)B �M����Mh0)�%������
�Z�̙���v�_Ht�� 6`�hghါ�MKj�����Q2�p�;"�t�r�t��ȸ���tq���$��3F7_��q\�aΕ�>�8��_���x9���.�N6M�MT�`81���Ek��A�2�Պ�/5y���%&�A�_  �M����3o�st�D�q}��Ύ�c��9pQt�7����"d>#�UnI����]�FF4S���F)i|�glA-_�1h�xy�&A���jt��b!mr@dm�<��*d�\��A��,C=�2��FQ��to�0��������~ˤ��Jk=/N�b�r�_ |��p�ͮӏ����  i�U�����z=KP�����`���۞�66���)��U+?O�15�������$x��a�UnNҶ�L�x�)�i�� 
S�\�A �� `Ǥ���F�!�ϩ
��:[�� �W���*������M��v?� ^��פS��(�n3����]�X�}��8�i�0���<����\O>t�۷Tc�4q}�O��c��@���ؚ�i�Hk���#}91w��؍�����E���������I�0���6ڡ8'}f�3�����I�~\�0��~�(���z�;���o�gʌ�O�#�4\dJ�4���I��3Rվ5�Xo���ZxB��W1k�t~��=��#d�Vl�Q�oE@�%Uh�ۄ�����!e����^�'�W�Jm.�%�C�@��<��hM�K}ǌ���=���.)��! 
3M����,��&���Z���cQ��՟57;U*1'\�K��%���؍��J<��7�7sW�I��/86�q[ۊ��0㜉���n��xF:ށan�XYM�pD ���x��i��tp�S[�$�)�M�k)#LP�G�J��-z9�KS�AY�`pB`C1�2���#0�@VMN�^��@:����{D���r�h��a����'`��Q�v�l��W�<�cz��� W�g�w��%i��D�4,�w�3_�S!0^�7�tpW�R��.�cn�
�af/Է���"q��"*2�oZ�V�ex�����ބ�=��|����v�9h���urv��ԧ(C6��/��Yqr �RY��������df�?�#���~�߰|�{׃=:�
Z2�F��y�O�6�Ӄ޶�WP�B�~��̘���e%e$T��bӡ��(2� �8���K���!f���"R�8	N9�.,fLx�H+�F�tRo�/�O��˾�m�QJnҠbG�S�p�oP����Tű�I�e��#����$�h�� �kɕ��p�c����::����A	�l_���wl��e���J�܇15�<�>�� �!���E��kz7A�ZɤD�k��2�&>��f���]XH��]��d�%O�
�L˵���6Mf�����cĵ�H\��~�î�5/�B˴�JL�0Ys\�k8�ǜ����Y!��`Ƨ"[���W�B8�ĉE�OLr3	+L�<����'�l�ٰ��|��J3]o- ۿA{?�pD��)�C��#U;A0�?5B����Ď�tJq_�,�c۷2����o()������ŉ"�H{���� ��UKy��3�'�Hpe'7;ICQO{���w_T���ǌD���S̽��j�jA0?��ϫ%�x��ճ@����x�{Y�@���F�7�����6{`;��ΠH�J���j�:5� x�x,sppjs��o�Pl0�.<�>ѭ���*���Ўr�86W�9	��Es�Yʼg����?���aS<�b(%�x����`�6Md�3�ihW���1F��O��8��;U�9�ŗ��P�r譢y���!�h~����<D�ː�"���^��������Y n��c�y �r�>�7I%�ēdw���&h�3Ϧ΅ڂ��!٪p���?��<�Zx��,�9�I�����;E�� �bγ8B �=�U2��a윜�z.�ZŁ[���ry+��L�2�����\��p�0��}�e47�^����Wū�����.��L���Q�j8Rj"w����Y�1]�B��W����ldEr�����gض�V��嫟�܌�MY܁�e|�➓M�BmK�G�/��ə�f���0vU���=�~�t��iY3��YF�u����D-��K16u(Z�?��j|	J�΂�2V��1Ն{��/����2&{�6߆��Ψ�EEN]�\�	��m@��l�*b@䭤V�ߗ敼g��d��b�:k��H��i�պ���s�-T��*�����M��.SF@�O%
����c���=��'P��U%?�|�/�w طñc5f*Q<Z�2
�	lG�>�]���ubM�A�7ٷI<�$����3���5�d�[�)���/��t�E��cPp�`q�F�EW��#D��>��w���{���4������� %^�Q������-�%�[��v�+1���J��~�\U�ݰ�)�NP
MTy�Ypw�z*=jy�r[z�k��V�.�7�*��^�/t_[q����_Y���}:���@抑�D)ˎ��PX�<���S�-�����K�&��JU�7A��J�d������p|���Paܕy�Pz�!�,1B�c!AA̝=7pH@!��U��0��$,W��Ԑp:����M���G1��,��_G�.�|�@Zg���t6/�m)������������BM�0�dS��$|/��-�����"� ����n�%������G訰�3�"2�	&�Z�/^x	�II\T��7�ڋ�0E�B����'��B��8g�����6m0'�A�|
vտ��gs5p��X�2z�>AC����޽��p��j
�%a��ͽ�� �J$F����I.H��x>�u�vWTݛ�IK��3nYp8��|�Z�cl�\�y��(����^b&	��/��A�1\N�IV�s�[sG�nI��LTz�J�H׫�=7�G#�^B1�:�lu�3o���L�&&^���V�<OlwIXAɐӘ��G|���k�J�k�N�[�j�۩�.��a_rk_�T ��D3�,����e�wY�Ur5���l�����c"�~��j�'E�FK�+Q������$*���OfJ8�Ҝ� ?g����bPJ��ܮ�o�
�Zf��� t>zp
V��v}x��kyTa �L\��L���@��0��un-8�i��'���c$J@{r��Yq�\L˙%�R���<{s���9y���f�-g�w/W$�cĝ�>1ƫz�t�]I��O�[����V�-�����Cn#��r�k���S�cW�gg��o~�L<��sc���f5�
��(��������ja��*g)���j_�㙓��	)�����V�����Z2&�����2a.O�!����=�����[�CdУ�W1
��F�wnҦaiW���f�l� ���)���pQ��N�z��i	=�ٜ�xzݾ�,��^���4�|M�������
�p_Y��/�W������1�4��_Fin6�?��$�Z�����A�XA�A�;RպU�0P=�ɉ/��{�n0PL��f��k-��γ���׸X���;KU����̊ ���"��NVܫ����0���p|sw�P�b2`�]JE�AY�Nb��* e?��i�knQ�߳=_>�^�M�
 l���&�rh���XOE �rv*�8:ٓ��Vq"�%Jс�*�Vd�A��l4�M���.JZſ8�74&*.6�J�G�@[�J��k��Fԛ��a��<>0el#J��c�܏1�.ԇ�i![[�kٖ=�j�T+�I�V��6݊��)�����V�Ui���۷*
�c7���9x�\mm7Xuk��;M# a��F���տJPx���4�F��F��C�O��0�"�#�P����q������:gb=܀��,��$��{�
J�)��۱��[����� �|�,"�:�ݥ�kl�
����#�bj���,�]M`�9 @`<���v���@X"6��)Ѻ�%�jR-�$�y���|��,�ŗ�[�[߽5��
��z�׿d~�C�\�0e�}f���-b2V2Ư�נ迤<B�m]%��̿A@�*F���
�gp�||С�K(T2R{����SKS���T֪Ϯ��w8�E���tH�?�I�p�ž���(�y˒������Oě<����3������[z�Bn��`�����E.�����W�,��\m��M}ď��u�c�M!���I���
/��9s߼��35PXjŅ��z�9�7Q(_o���O�I"�}�|ȏ��b8-j��uk0����{I�8�H���~�r6����	lH|zB�k�\�5����xrIƓq�	8}�!fwh����,����O�Fm�}���KŇ��ʯ.CPf`���BuKc ����8])���9h-�s�Z]��Ƴ1 {e��8�ED+,��D���jC��I��G�}j��
���׾=Tj�k1���G�fz�m�`���q-p�:�V�[5O)��T���y�1�b�x�� g�dQ(�3�7��3��R�Di%���:Z!g ���,��r{�� ���6zK�D %瓇Nۏ�S�/T<ժy��:�l?�&;q�ˤ���0yk���A�W9+�l�����f�Ӷ'��e�Gƾ儫���]���@�'�{�+Oρ���cǶ3Vks6]l�p�:	�F9hxX%)�Z����B����-�!!�S�]kY�%�K�1P��I$�ΨvΈ�(�c�lyQ�PN\iL�ݬ!8P��A@8�ߒ,���c�@�W��啀㻢�W�~�|t�B0�a �Z�ZpZ�}V��̰ �x(�9Y�7�>ف�g��Q�/?鏀�m�����PQҼ�-���I	���~c��A�Ї�4�w�pk%Eٷ>��ô���bԳ8�clz���$9���d����%��(7���Kb���&�{((MZ�6��u%d��R"w$�s*����!a�9H}��_c��ϼt�KcRj���6���9��R7��(��W�[�=�y[Ի�i$`�hC�,�1?�6^��Z��ԇ�Ge����؊�K����'%���Y֔��^#�����tU��t�Ik; ��Sl�Rs�Q����#S�u���v	�l��Y��Ǩ�rڣ\��b�睤?����̌T	��+��=�j\*Uv��}�P�?
�:�;���>i�r6�c[/���m#e�*v�)�j�6>��	ҭ����էҌ %��x��1V�K�s�x�Apr��_B������>W���CІ���3�.�b�{с��ۏƿ|�_��O����5�㡉�7#>��+��(,0ݒ�Dt���t�����(T�D�M��H\�;?C�|C���pg�Dh��p43�Eu�x��B�C� �1kz��ڹ�S,�*��q����v�<�γ!~�Ub�6�HE������u{`���lf�������������@u��_�]�2�q�#�E��"��������pQ����e�/+��rc�+Զ�uӫF\��*��H�����T��*��2&��/��ђ�j8³	��CK�<��#}a���>��_�)��-��x=]�3Z��F��<4�&Ū�r��T���p��30�.��2�W0�<����3I�<��)���!`�nk�={#}8g�r�܈\��A���'1�|h����������#�˞+xznǋ5Y���k^d�rfE/�:�V>�.-���5�����#EQ��,�ħ!޺dw����ulf+:������ec!�o X�/��~%"IpB������Mnq�M����g�=冚M���iy{O����w�f�j�c�7�ŧ��X����T���@�:<#d�T�=:�c�����YԻr����9�u�5Q��?t�V�o7|ڣ*�h���nM�R���Й{��7ֲ�2�פ�0�Q(N���Z}C��<�1�G��3��
��͏�7A"z6T��e��?�-~_j9�����u�.�^1@��L׽ |�%��86���";4�%s�`�����;0�m��$���4G�t�N�Q��]�d�
�i�����3V/�z�F/^���4([���h�F䎺�Ҹѩ.8;!S��zh�0S��,$�>o�>��-e����٭^�����k��s��޴�
�9�ٝ/O��xؑ�,4��LD]�����o���G�hݭ�u��-ń󬻩�H�I���K}����ܖl�*p��4��@�Nj��A��7K�K7a M!������{U�����u/��H�}�e�߃�X9dě:����w��W��!"H�Xνj.rO�X�H�<�7�8��@D<J�k�:�.�+yw�]�]$�5�M:)�?\�����\İb��
�d���e2�I��;B�c5����:�1�{����~s_�	�ڭ5��D��fP��&;��80`��)��Y��B��<e�)QP���khV�j�PL˳$D(t�ַ-�#KL�V����+[�����
b�������u�ں���t�pf�^�u�P�+0�?h<�o�E),���\H�"�$�� ��f�0A8��{��@����4]�D,M(KG�:5[�W̩��q��ǩӤ�� [�{Vrp�Y�vB�n�s�~��v���g�FJ�,��G�D��r��~�]r�[3y��Β`֦ͮ뜃�ڲ��ښ�%��Q΋r]�o�$f���C�?��������M��]$�V�;��be]�O�UR�Fm`�!{��ސ$Q�-A:�Xw_����y���^�2+4��lu����[Ī�6�R����֧�����M��T�e���.� �#�՜��7��O��R�����ޯ(�'�����e?���xa�55SL�n����x���poF����h0�p�����5$���!�.m�"��0�J2-��&��'��ҷrE�h(XlxVHYEB    7d55    1450弥�\M�Yg��K*��7%����q	�#k f7�`�3��G�*���[��O�u=Łt���
D=�R'��s��˲�qކ:��F:����s)�<��߶|6`r�G���=��0�N���G�
7ϐ�ܧ�Dg��f���O�J���jjNޘ�� ����8jl8q�h��9�,N����G��iU	�AJ�I,Ʌ�D�:�D1�FG�3�pF/�S�`Q4�� (��_����w���
*��XjS��T�����~+��u��0��r��h������0zP.O ]J�ΑR�w5�r�'p M7�8�.W*���[O8��u���_T�W�2ڃ�f�_M���sK%�E��@"�:G�U�5Y/~%���/��M+>\���Ŗdv�Xq.G�����m7Z]��x��ң�� �ź��C��iup}��4T7�~�0�:�����2�����̢��e���%�u�r�`�2w)w,�=H���r�O�+җ4���B�S�j��1Dkq�q��S�s��Bu�����e6l	y��C ]��B}�zh\$���Q�"�==�v�}E)ä�z4�W����y���enA�~n�>B��ʦ��8H��f-�ſU�#:��=|i��>�K��8)�3��!jo��3����Ucus��&
�;�Jt��:�� �PkqEQ���*�M�u�f�@�[FE�;/��Q�6��1��z����$𔪜�e@G�*V}k�!�ӡ�H�E0C��Z�$��h�y>�K�9�@Y��&�Ǣ�{�F���%Pjț�o#�k�1s>�iR̈́��y����@9 N)��C� ��5�qܼ�������1���6�����H�:�G���ٶ�*wg�=���3�ߘ���>�y�x|����ǃp��Jȅ�%��ϕb̏�]��\!|���h��5�]c(�v|�Qs_�xp��p�i4���u����F�<��opU��g�<�9.\SM����$�"7W/���oTp7���,Zx/�︚�c{3�y��6�M�4�Yw�F5F����*=�byD?��EQ�Uw\<�\Z�x����r	�6//�Tg�d�H���_늰aآ�a����{3����t1܇��l��ĕ���P������v��p�Y��L�<-(V�B�԰��������W�s��@	��J�{�me�`�/�F�y=����׶�B걏��#��t�C�׿���7vW(~V�����nY��>���;ɣ���o6�	���!e=(��C�?�n����ߗc����A���e��,�C�4����e�ڎ��Ml�fᐪ�e�g�h<.��K����6!��ʯ�4���I�1�|<�Ʌ*��'�"��F�Y�Jϕ5��v�/�)(����.*�Wd��[w��w�$��{%��.Oj�fGj��y�`b�.��F>�(>V�F��m�w_Zofɥ�;��х��	�O�y�^��r���?��:��j�~ł�=���sՈM�=��ۆ�$���SA$EkʘA�e\�� %XG�Ĭ���٨Z�8̩cz�M9���	�eZ!gں����!}�['��J�Ϩo��פVx�����(3�e@��j�S�5j�LAv�R������,��L�#(E���A�����_\}��f���D������a����I��x�j���j����N<�#75������wV�X?� �����Â��O7B��Ɨ�[	���G7\�b>�|\+=�F��zT���t�:]���X�%=�e� A��~������V1sT��_P�Ǡ5�HF0�0�6�����MɅW�|�;X1hA/ۡ�ee�5����JH�� �98��.u0+�G;(QE��i�Bm=�V�8�b0u�`ړ�v1���u{�4���	m���N�&$����Z��� K�k}��X;�x�ݤ�V^��3��G!}��[[w���JJ����HN��K�L��3_�	�%�p���^F�">N螣�
�ĵ-�bx��9�k��r������X�W;!�N������æ�7^��Gr���/��'�brH�, �'K��
K��r�mϸ@;TS�8�7~�#��G�6���BW2VQ3������� �K�ɦ��X��$I17���!���lSx��u��I�9�ʔg~B��c�7[L�>e�4s�����[��.��gv�`�,x.s%��0����j�b������ȗ�!�E�i�'5e��qC�p4ﳩ���QiI�!UY�G��y\�de���.�cS^�^�b�q����g������ӿ��U�J��M� �#�߭�$��usu*����o���s�B����`�J���9�CJ�� ��3�o��@ĒX�\6�����'�/?a5���d��sS_�j�u\�q'b�)@�R�v���;�� V�����>pm�]59��8�ӫ��YN*�D|�Z��ܾ�`�wQ"]����o��,����Y��0A��_�@\X#�>`K���œj��)eo�� �Ɔ�@���0��ϙ�A�nʷḠ�k�a��k2~!�,���մo����3�H�2E2��x|���zi�۰D�7����������f�Y���)���-�ES��\4M�A���g�T��vf�#V����H��e�Jp����IYE�"�DW��b�H�4N[��Ng�܁�0�Fu�7�1e�t�p�Ń�JL�⊪�Ѝ�Y�M@cFQ�C���?��^71�F 4�C?��͙c��5q)
E�}[���*�����9��7�fż���r�A�N�.�"�5�6�k-�jM�N-�"��|@T���qv,���X��a��Io��Jl�y%]r]��s�{����ʡ�4��m��F�ʷf�4���c)��Yq�=�peh8 g���m}Rb��P�����Y�G˛��ޣ?&�G]��G��h��
<6�j#�ZtzW*1�g^��DG�%�eT��g�|��E
�V&(�D7ۙ�
!J��9N&�*a����K��9�u`&q�:��XN �3E.�eϱ�
�����i]pt'�Mu�$����A ~�-bH���a��w_AѴp��б�.��%=fs�b-Hݎ̲�茄��:�_;��X��w�-�J>��D\��{]t_:A�$��k�FgA����f@����*�P��!T���V�Z�d�kє\��^)��[��gA��/@�����=�좠��~��7�7W��
xzZr��r�+��4+��wc��� ��wC�m�A[�0�C�=.�{*W�Y?�0FI����3��0�,��69������l�w8E\��> �[:�J)S���S�C�Ծ�K]�}�l�t��j�|&������$��(dPd���1��O��C_���|F��[��rn\��1:�i��-�LAG��x��5yh��sG���l�1v����$�=ϐ=��k<ZuN|��_�7<��J�Y�,�36|��Ɉdl������u�,@�xp5�RN):r��?�ib��n<���cp��aj�T\��������擼�!	���2~�� �&n�z4����Vچ�%��4���T|�N��̠�r�=�9�G��
6�>�V�#���f�uN�Y{�i�0�E���wI����b��/��A�ҭ�?�7~�`;�]ׯ�KC�D޾�u��Y��6��3\r+�������qvzDpwIwc�p�A[-�$ M�c�����wJ_U�mdLkS�9�:ݢ�FʝPʦ�����,���h�Vh�X�
Va�{ğ��w3h�����f��K#ׅϞ1�7iG	>j��$��z� ���pC�+�&��|�nu�����nuf���Y�
~�dl7�	:�B"��m+@�N|���Zƭ���{�W�:6�Y0��."/4ewX���j�%5�M��u��z�(�a 
[��=�K�Oz�yS��
�C��#=#E<�
<4���]��Z���.�>E�k�z
}�N	��$���8r������*��B�k��ȇ�m�
�����
�6eJ"�z8���#d���W8�*�%�@�@H��ߕNQ���n}�S�`��~���ճ>�@*�*/.i�ޚ��W�ME��qd).�/r���X����E��+�,+1cS���w_t�]�|�{6�g!�9 \�nOU��A�)@���rF�N⡈��xd���*b�n�Q[�i2P_=�It9d�.�?�9L�j��{=�W���E{W�T�Lv��%hE���NN��v�^m��tE�oD� �	�CYpO�妕�+�/�e���ʫX���z�|d�~TɰF�0�=ޠaI��:���QA�횊��I3�5��.�+Z	j��	�05合D�{��Qa��>���&C��#�d�B#)����c�F���<�bDG����FHD"t�Kċ��lx�J�w�;��\赎��ܓz\���M8B\�o2��ǩ�cC�W�s�B�
`�U[��|#��?f6����˪u��J��'�]|=�-��HIv.iXg���[1�0ٰג�{;��p�#�M�KY{��~��sÔ�H�V#�kd+�HmJЭ%?.�	�¹��(~%�i/���u�+���ٹ�@�7{$�c^�᧺��0i�Bm�B@���.݇��&��&B���m�_v���Gяx�IzޓT�&��)����.J�vn]h>���n��N���Ĝ�.t�i��\mD}6����Ux�����i�7��J�Te�EeuXg�,�$�m�Y+�T��ؖ��q�+�	<T��%�45�,��f��!exb?��su�Mw�0��
�Ln 8b`��o��FEOG:����X�� ,�Μ�wH0=}F�Ȇ���>�g8j�s+~~�=^�%ks�\~m����߾�p�7������x�U�����#��a�ˢX1/=餇��@�%ٝ[��<P[jJ
:Tçg��Ϯ/_�y`F��H`��l@k��$�
�*��pUe*Q����4\�פ)l�\�v��[+�SZAJ��i�lHߩ�E���������`��$�7�	,.�wz�DW~����Z���#��;�<U�l��YO�zVy��=To���Fq�[B�XT��5P�S�G�+��>(ܟQ	���pp�ib�ԍ