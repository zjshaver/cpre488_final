XlxV64EB    1852     800���9^O�UM���bz�ߴ�r5.e��/�u :���ퟍ��Ʒ@k�Y*�3��K>G�lk�K�6	~�\�J��!�b�s��7���$N��N%�5�x�X�J\��b�[�l��/#��K��{����ꀿ��2�.<���A�/m����^	>�=b?z���P8�3w�ys'J����_^�wҘ��z$g�6d��
���qG�����`J@���C?��]�E���h�ꧩ��r��}����J��}��kA��$6��E�4��h��J�ʄ��DK	@ڎ
Ԧ�B�0w%P�d�o�Re�~���;�&ͦ�g��a|��(���w�!	��Cf5��-���-ݙa��S�xV�\�#�}4�T$S)�&��8�3W
���i#_� ��p�0B�W�lG���]�eD0�ɍL�IK?yJ[�=�h��������%L\��Td|���2��T%�IC�f�hUnD;23��
�2_�7�)󔍾�b�Iw�#v2��E���M;��BQ(��23�7p�f]r��F�xw�՛bc�<���K�C� �2�IJvKy�g���\���!�dk�}�*Ң����Q����0H��_n �-��ώ�<��Ѭh��[y�����ahv�=�͔5��`�8�i��'/g}>��J�ќo��\�!e/�23�m$�����������D�H�
�
�T���s^T^Ηq�@Ղ��1�,w�|�) d�DJ�)���n.�BjK	[v8�`��A&C_�3-�:T �:�p�B]�d)[�Nr��Q?�:�U�;c�<t��N$��Kx��L`�ȁ���'r�$��0j��_�F޳�4rP;�ņ�7�P��5��˦ Ȑ����Q�@<�i�+u��W#�B�/;�8�7�ʅ��DW�1�2����J^�� kL�L�Q�V�����O\��Z��I��� 6�X�a�����LY���Vm���o���Ps��K0�;a(L�s����%v?W��*O���A8D�� ��a\�Is����sDAm���y�}c��l|	PI|�0�A�gP��b<vV��%�b��[�5$�5z뺪"V��\k��Y�,]�O���r��OW����9v�ߤ� ��(�Uևdx㖻k��S��M?���T��p�f�D��c?jRyu�XmBY��mml�X;�����J]-�6�І6s����/��FZĶ��e,�oc����:`@��e���ݟ���rG�'��s���L��F�-(�>�~<�ˀ�&fS8��PNF �&r<��4��������6���<���
3�6
���;�9^9��|	ޅ2V����v��y���W�#�tO�v�i��:�\CL��"�w(�i@�F��d�����z;^o��U>��E���|�6�H�x������J_·Aҟ��:+�lY`�E�HUoLR�����8x�������X��abB��#����2�:z���'E��v���& P�J�f<�����U�)a�>�(1G�����7G���>E��WqO�k���y�$)�G�Nym2�-�Ma�~6:]x�{�ܽDh^d|��7{E��y"p�L7P3i!Ď,V̬��=�AH-Df?���������c�l�����򚦧�D���ʠ������}�:�~h��QE'��m��.X���l�J��os[�����0�&&L2 \�o�GQ���:��:�����̘��A����x�,�� ������V�����+����s���뿞m��:�x|�3�H=���)�w~�\,�U�!�.�^,�;k��xt
Wf0�'�7X���8lԁ���P��0�[P2@��F5ۄ��*� ����J.�4ʳ�&,T���aV�G��!�軶��<K!l�oۍq^`�혤�����+܋�(u��~V�>��âEv8��s�h�?�-6!�` ����|���?m9Lv�i����r<��4�l�m��RY��5s��{*ӎ