XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������N��,��$;�X��1�E²0�Bc5-V��F�[�8l8w��E���V��KUh6\�����B���P�푪�|����g�NGB"����"Ѿ���p��A=�oy���`˦wwUB�G�QO	�����	B3�{l��;�gצ���������F]��u�=K#q�=����&�9NB8؍�Wp��q]��毦�?��Z,i� ���N�f�%(��%�.�=n�����?��}y�L�.Y���.���H����M�w��&�9Ѱ�?�g�V?Oc�
Z�@ud���]�R�&��ߞ��� ��4*�mS�9P?M�Qc9�h��i��W.(�,Ɓ8��9m<j�8���ґR.R �RT������,�99�1�zI�`�(������M����>���c���Z�[��2��>�0����Fx����\��L.i���@�?Uj�-',���Ҋ/�'��&�R=�I�	]���c5g���W��Zi!�%�.a�.U0�Oe�M�'�\x����i�L�X1�( )�С�ƴ]�{��-���t���R�,>��j�w\���2�=�:�-�Z ɺ2$����4P���fi�1����Zp}d���!F0$��]�{��;�d����H�b���B�K �ސ��G�*��Zͼ �T�M綀������5[�߮|�Åb<oM�ͭ������T�8'���:'4q��������I�G��œ)4P���1f�`�h(6hE�ߏ[�����k�5�XlxVHYEB    3a46    1050��m�N�R��µ���Y��KBl�Y�F-Bt�:���6��㴯���ܻW����O-k���Iοc�և	�X\|<25��&	|Gy�<6��z}�D�F֥.�!o|���� د��0�S�T��m�I�eOx�ޕs�g��$J�Z�<=�����������>�&A<��9�)���&Z��Y2�6d���Q`��Y�A�<�3�|���}�l�M���%�9�{�6��Y0v�s1a}�R�@w�.Ō%
�Ӈd}�B��ؽZ����L��/��2@�fct��&-��o�C�\~ଐL�%��v�3��X1[p ��.:--�?���Fw`��X`���DAύnSg�f D����h�)q�����@���JJƃʕ�>�Ĉ�1[�r/�AH:��@�N�bD�HDOCԗk���AZ�7�H�[�9c���pl��Xצi�q� bҍ[���[]�U�|����ӭ=�������V��i]���ARht� ?��N>�5��m��`,�1�_���:ܻ{�UN�z��}��7ؠ�S�QZִM���� ��M4]*iէ����v�J@w�*�0���/wZ�PȫSN(�a6�X5�8Q�u�s���:1y�>�f���Ѯ���
1:1�#�[�r��YI]��dd1����Ťz�ZC��|�dXt��h�*��`>]�Ԗ�{`.2wk>�v����lh��3����(,Ӊ�J���W����ow��-dA�����7h��9:Ħ�G��H<H�[�`���/�`�Q�GHb�����>�h����c��[E���@H�>�$^�Ad>��C�۠b��%�y��v��s���!<�ބ���ڿ�Z g���[���Q-�ڣŸ\աq��Q�ϐ�@�%���h��F���j�K=�é��q�]��MZ�-T���V�K3m�j֓ҶU �L?�DAs����bv��C���X]Q���[����D�1?�5�ܺY���`A\.�WSB���Oq^*M�x��)��M��GH#�@�:����ץx��ᴁ�a]�T�	�������	���f�j��h5z�)�8b��	��e��&����� �{�18Y���,^Ϣ\J�u�W�r�������֔$;2�e~�J��Gg}NA���� K����\%`�O˨��(��ӳ�H�L
�z������S)Ǻ���wpt��Ec�D�\ʁ3���}� �;�Jy5n��Ү}�����v��MO�9��9��9���#Vͭ^i)��:r�g+�H��:�p8��+dM����{n1���^�vƾ|���DD�"d�(^Eۃʅ��ۖ�2ԁ4��%�n=�e��8ꈗNj��oe�f��.o.�j.�*E���'8��Z��*U�PP�R��`t�6���ҵ4T���,vXh<��e�V��*��H��!�Cu�k���;���;���r����|q�1O���Y�並��Ɠ�"�'T :
Zƌ�äe���y,C*�6�c�#��뚟X8�~;)[��?m�\X�r˓J��N;(�����
��@e��|h���9��ҜQÝt�$��y� � �C�bs����}PS�`���e��7����t�%��4���ݦ��tF*ԓ����ٷ@ ��J6�Eʵ�$	�~�ꐭddM�1��e oN�8�"$ +TF)��9����3�M���&��G�OÌ�HLt(�5�h�Y�Ux �co��c�� ��6�-���;@Q�����)-(������>�CW4�|q��[^WE#r�&9����l;�_���h��gY@9�yZB�)=]]{�D���#�%���eo�S��ɺ���a�7Cz��`�}ŘN�-*��,����i�uK>.�y�%��G�jr�j?~�%��j2��B���<.���,��o��"'�^w�{1`����s��S ��[M@gQ&��+�w�z���nܖ��?�X ��Tȴ:�T+7�;b�V~W`<���?_�y�}�ז=��|��2�����3
�&��m���K�U�L�o����~�4��4sH�3���r�2m�d>�CF�G�n�7l�ƣ� =��_��~}��ha
�tɞI�lf��-N�#&���LZGTH��0$,S������ӿ�Ȏ��S7Hfs_�E��um�_M~��j��������MNJ]��L%�/����;:!�H��)e	g�ܐ�u���<���2Nw���z���;���(X\v���mX�E���2�WCx��Ѽ98�R�>ˮ\�Y�2��)�����"a�F�L���T-��
�e��>#�'�VI�]o�m.@e�#��V���j�g�A#�P��;���h@:��\�؊F�S��#� HI��uhW���
<Ǳ���c�q�c�P��~qD�*�VNE]�&\�vr}ەYj�Q�N�y��R��0o�_�y3���ʞy"� 2.e
(�@A*:8�~�AP"s4H2�1�o�c�A�`ܣ�d�cԏ�$�X_c����͒�دB(�O�S��Cɱhv<#�9��e@Ҧ钜@ݗT�eZ�dv����� v��b:ze��r�h���~e�Lz���Ʊ�I���s�S_>�Y���i��ɔu:?[�6�#�t�r/Q1e���ϼ��V�E��Ȟ��	�����S��C����J��pD0x���a�\����ӿ^�Sl/v��j1�5��50!7���}��m���eD��x��s�-�E��Wg�N���Q 4���!n1F�s*.|I����򗆤f��E_�ko�|�������ʨ�h�0(�]��`E�lAXi.��%��O$Lg�wC�9j�#�\�p�+/�\�Y���if�jaW9�R��X([�ͯ�Tih�c����� �j����L�����3��%_�4j3��eimt�`M�NY�me��e#ɂ����)pA1k�8�!ט��k�g�LY]�����T����^��M���{
����>l�ɥiƚf�T�6�3�(�1;��Am��1��`"��5��jyDTx��0���TӃ����98\�d�Hq���M�8�zif�[��:'�@��њ����y#��(v��u��N����s�+�a��O�-�W�#�3�x�Q�<��	t����4o��d3&ɎF�1k��#Ejl@@zSR��XF��-�h����vS����@|���M���y��=s��.z���1�B��k;��@���:?�R ��I���XƆ,1W7J~��=�Ρ����6���6���?h�8R�M�����එՌ�E(��o�b��	-D�odf���ܑ#��[�~�%���Msg*
.�[��k������z�j��� ������6]!�鰀��Wa�l=4;"r6 ��%�����WPO�a�����C�$F���ю�;�w�V�0pd��w1غF��ADI,BSu�;���	u�&�k/�0H�
9,u�f�L#=�0Ͱ4�*�|4�#J	�4�~��}Zl��0j��ch̑�*c��}]����u�e���#�������D� ,�uGK�5���n�C���;^�:Lqx� �_��*&n��`%Qq��Q]vʮ��ם7��*��q��m����SX�NnA@���U_m�cN��
�l��M��/}	h�`����d�Uk�@�S'=��X����`�%
��/J'd'��3h�}��u���\���rm΅'�>ygĮAȡ^4����o�?+�٤��~�u�%��)��Ǻze���I��ז��@�-x��ݎ0��P��%�j��&2�[_%�����4�h^p9,��D��x�"�%�?U�j�gǚv�oL�f4K-�����٢�"�&f������V} H j�ߦ�4�~��V�^6 ~�dU,�XO>�u>k*�9���☆�R��)FO!v�/��oI� ����ޔ��JUz{9���R���$j��`�a 9}0�NM���7<Xg���|=tk��[��z����EZ ��J RF��U�Y����§�ۯ-߆b�zM7f�G�c����/U�쪙��X�m)1R;�nN��.[!|��'���U,mύ\�}�>�?�Tc�L+*