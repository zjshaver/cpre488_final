XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������j�k�B�DC�w�7F��1�}�nqM�QyL\}�X�m\3`ȑ��{�f�^h=S�|�>�C�l��$�y�1��+*���U� �r_f�	
c�*X��6����>p[�۟L~���$Uކ�>Ųv�M�!��.Е{�mX���������d��d� ���zT�Ư)x+o����)�as���B�Y��u�'�kS�k�G+�t���!Rޢg��L
JQ�U �Ϊr=�S��^^1��q�;�1S9��)\�i�'���7=�Y�jgW}�p�
�����P:���yʳ씣����Ã|>�mn=�URHJ\i��>��/5�Ɲ�V�ahEU�_@ܝF�Nj@V\\1�=�rH��'����z+���>���so��v��pݦj��P�r���U� e3҈�*�����|B��Q���aba5�U�${Ҥ�����}���}ܰ�>'rN��H�究/�p��.��T�7e�`!x���/<�j��^��!.��~�Z��E|~�Œ�>�p-j�sҚ�Gv���P3Yz��5�٪)��<d�!���1�d��Jsqc6o9�V�!Oaū��x��a��� �r��侴n��d�塻l��x��qe�^H�H ��s.R�<���ҀO�x��($�v��w��;s�(����2#�mp��& �������"���P�\邐VK���K����G������vC��)(����i�hR�[{W�H��#���x�~p.�]��Yǲ�?xV�8��c򮔭�*��<IP�XlxVHYEB    1e3a     a20�D5�feenB�z}U-wf�Mu]��<�W�y�DL)�5?��g�a̒�]������1M���w�B�N�v�g
��,,�U���ZB!s���T���+�����,s�x:�lܩJ�)��a� �ܶF������Ë�v��O��)	:y������g��h����<7��rECG)���zH��vmG�����^���p�6����h:jjJ{��[���L��n�����1Q�!G��E�Z���a6@��x�������S��1�>���^�g�Y����q�¹]�x� �Ae�֯7.�.�pxQƥ�ˊށ�.2���P�L�E?6;�@�H�]3�����x����#���
+�Y���?S�ŝ�?�R�Ժ7�⫶�7|[��"���ɇ%�oP��/C��ZXDIk.���4�����yv���������JS�Q��g;�GR43�`���
U� ����c�*W2�Z���)D<��u���zc<Q.�?�)��J��ʥ��'�W;f�		'�KY.���JI��7�� Ge��'*vs��k}A\*Yc�enY&Z��:�cr�+�����G�����\������wȟ�U����%ƙ�,��+�o���d�Ռ��ђ*�<MD(��%�p�v	���VQ#�i�H���Hu@�T���bJ�G#�;ŊA�V�¶�Ge��t�^,X�n�6rl)#�bkc�?9E����J ��i��ڀ��Hh�3�3;�2�_�F�H-&���W\+}�-�Y��$:��r�'�"B8�^�:��
�XQ�����
��~CM��<^��2Þ�����[�7�:�0j�~e԰*�̶�����'���0����JA�~�1D����~�	C�7+�&�P�LJ/�B���ʵ�_��D]V<��osͷ��:�h�N�fM����Q5�З�G���9(BKv������?F��)7���`���<ff�]鰰�?��V�?̣�YQ
��C���$�&�{P���0p��/��Z,G��DJK�5��Sx�[M�"����3�V���es���/1���}��E�	�u�i%���[��j���)��I�8��g�P��ǜ�b�q(/�ף
|W\�G4d-6�>��й����ԝ3�T�J�£`�7%%��3�8�A�k��#J���Z��|U#z'�7�//�[�ו4����$��.a�D��@��?�!�q�����7l}(��.p�ǃ �械v8�'��eT	27g$����[!��(��g���^T2��df��ua����D���T�t��dl�B�m�uԖaG����j��W�K H5�"	eg�\�l�k��㜦$u�{�`�g�ϑ#�%�%ʋ�ʉ���n����e���&1����"�~��/n�-:��C���A��葻��qj����:&�䱲.F��o�mwa�h��np���]{�K��:� �]ص���q��2D{���]`Pu��Y�v/�[<�5:pC���a�x��0�>�*�����M��
,�[��y��ϑk��^ez^�'`�^�U��d����͞�s;��Y"xPp�;�ϭ�c���k�h�* �7S����W����6j�Z�Y����sxbQfj�O�B8�V��q0�@�>$�
��!�-U��L4����a������އ�����2	�����6��QC�f)BOc����c�"����'�\(��Uz�~%2��� �er�鴠T���e�-����}����ާ%v��\���0AE���d�?����У�7�3��5��>�Va�g�i������ wDJR��k�����r���Ch�3��Ͱ}B~O!9�@�_	S$����5�ui�=�8���
A�����-gO��0�/S��g�^�R�6�ȅ�J�t�=��wh��M�\L�V^�jr�~1O�fQ����M�q���c�Rr�B;?ߪА�ޣ��uE�W�L9�7�������+uU�<�m���&�_���`�kX���7���pK<�1�j�������;lS����GքãO����(<��J%�>�m�M�_��N$W�1�r��a���^ͤ��@�g�52C�L�}U�ed�|^�
$�0:�̈́��F��3��ǡ,���)�\�	�&-�;�`�a����
��F��9�J�����k���
�&h��T%���nR���U��c��2&��ㅓ^qQpp8�]B�24휯a\�3B�	�(�,�QgV�N�;ٜ�y�V\t)o:6'z]��21�Hs$PF�)�] ���oSoa�-(5��J�)+fBٖT��+T����|i�$�����1d�v-}�mD��&�k$fi^IJ�_������}����r:�G���$�zR=,wr����qY%��(�$���zZD޽о3r!�Bp�_qШ�HcFV����NЅ)�!¾�k���Q��+,i�d�������g�-���� #n�.�W�qV�.�-i�O/S�q���\�]-28��a��5��F�O|�}����� w�{��9y�H+���Ʀ�um�zZ�Up�]��