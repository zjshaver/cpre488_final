XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��V��J��}��YaK�P��2��*rs9�ĭ����X��𳗮5�T�'�!�,C��i�4�C{B��<Aȶ��Ț������J�l.���=���,���cll�Ξ3-�9z�[��9�w�V� no�i팺y�1�K�#Z�Y�k�������˓�W����e䃈`:]@�2�\͓��@X}j)�'���!���i������ˡ-���G�t�g�/kג�/��
βb�z߆u"'UMd>�0c�07���#_��-�^G�
��������^�c����ѓSm�u��G-2r{�D���dPk�.*�!��q��x\��I�P��Xmg�~R�V���VjE�ukT����}>K���l���O*������	�G�y��y��`��?�Bi�ӈ�Q+p�Uv�*��.1e!"o`��x���c��°^�:'>ie�"K�����o�.D�B�J٨��Np��9��t�������t-W�������vV�Ɩw[��R�ۡK2���V��A��F��]�74��K�?y�V�1&^�{Cx�gq����w�����Zت��Υ�e���Yn*��Z1�aj'r��yVd]0����L�o V_���slq���w�)�v_xC��fb��i2�ꅚD_���4a���Z1����Ak�� 2�엋�8� K߸g:ޡZ�~ �����6���^��T�@4�h��y^?��x�X>�M�����Ϩ�r�D����k����)���c�ܚ������Jf���9������:XlxVHYEB    5224    1740{��Dx
�#
#���-�؟�*������ܳ~�f>g:v\MN�����������x�~�����0,�"2�����]V,KM�%�P�	T;�|W?Ĺ'��g��N�T}���Ei�%�DܓpS���~��	o*�Ϙ+�g�&肂뒄/N�ܧ��IQ�U=O�J	9"P6QD�\�
��&�Ԗ�����0^t�G�p0OV���[��\,r9�!�#��,�(�'��5�6�,�����Ē/7��B����~O[>V�8d���aL�U��
�EB�We�݇�	l6s_ڪu*K(�e�S�x]�ժ�߆x.���X�WY�>���9A���j� �~0i!x��[0��d������I�Ж�x�z�;|�@β�FM1ve�vJK:�n�%�z?�#�6(^)��lB;���cC�J��f��d�Џ9{�K;�Ap�L(3P��M�I��,Ê!L��y�K̖��o���E�)���#ޑ�3R��a�{,o�N�����b����"�&�iC��sM�� a&h'��B�Gm%�2��A���h*�ǯ�E'.��r���|���٢q��}-r�x������c$��5)��#맜������۵�I\��K�<�ݦ���$uB�;�)jx�$3�\�(+�j�Y�JY�؏/"U��m�D#J:&������o����0(9SʡC�I8kQ@��j3�~f����K��	"z���
YI彍6PQ�'/ex¿}|I���	/�H�@A��	Ӕ�o��g��ڴ�S����Ln-�8h����n���B��*�E�d#�"�����&����w��F�}v�m���dڦ�n���˫u��z4E�Q������Ms3���v��iwR�����(0��~�$��&W�	ǖ���uζ@�׷��kH�N~&���X�wjV���&^���(7-�����NxR�"�����2�7�:�x�ί�֤x�#���N�rk�B�N�0u���9�D�'�Z�U��Ԧ����>eo��+��j^�@få9�x�nL���16E�Y��a1���`fг1Q0�������i���u=|h�i�ʧ�y��D�{�v=yܖ8ZĦ>���t��>�Cw���(tY=efyg�$�R�b?
yGL�@t����������I���_g���2�昽՗,�Ms��OlM��y�Hy
5X�>h����>!���D�;j���a��Ѻ)"7O
Θ/�ux��X}LK
�vپ�$�X�m�t�s���n~-��e�l� �D� �t���m
r���I��{q�`��k�A`F�Ż,]�pʬ�9t��
�V���8U�����ԙ�(���b���/�2���l�zW�핊t��a�D#�= ɂ6��yH��3��.�YwF���:��]���#c��̗��~�&��%Gc;|X���@T�P8�iji_�#0ʣ"��A����'*1|@���)�{#�����Ө�Z)b��qٽ�K�m��y�D��c��[t��,WW暴�`�!Ӝ#|A(A�13�w^��^����]�rS�a�F�6�Ï�w�e3��~%��2�秒���(��S�+ #�ځgd��!���qf�r��'Y�YO�C;ٻO��a�� �{����KA��d���`�hx8� ��5�!߆|ˠ�����ND*Df {\[�����x˫7��k�=V�t�HK����t	4��g� d�(�c/X����;��!���J<[&h�R�{0����(l�%et5<�7���F�T6p���Y2��U�uq�Q���Ӫa��)�*T5��z��"����������Ԇ5�qf�>��bѬ5�&���Pp��������W�T�݀-pع�E���.9.d�� t���ৡ��M�f����ձ]�������"W`\%��l��u�Y�MY[��v���KA1����Nx�E�b��KS��n�«�%̎�"ٿ ޿���ݶ���n�9��ۢ�,sP���T2����j3���:�Ӂ�KFH����/��#��xA�%D/k�kN��d =�Q�`����FCqe��c����@
���-����ݏh����3�OtF��u:�7��0S0�N�{������,�3��4��M^�|^�-m��ehs	U�d._݄��fz��+��h��*���	4�����U�y��~�qo��`z��:�z�-�d䰮��w���3���,̫3Qu��3�)5s(�N; �n���I���f�H�pBr#M}�Ef��I3�P�и��3	�V��L ���v���y�h�g(�9u��ۗ�ff�"EY!U8���G	@����Q;[�Nt;�U�0�x�Z�x��<��Z3n��/p��D@(9IyK��0�!e�GpB�w�l��A`3��WyF���6�fF��^�E�s��
K�(������"Ɗ�iT&"i�Ֆ'U|��qw���v���T�Vs�p�@پٺ1�S��@s;����j�T�yߎA&��%o�����<��I��1Th�x�z�1�h�1~���P��=��=@j�;Dy�j&����iB��;��$L�Y.�fՏ����w|�A��=��U�@h��tbgF�߭���w�K�5ƅ��F��fn5�]��Xo�?*SJ���C�m4b{Z���c �λˇL��H,�?�v��|���G��I��^�j�.����0'C:���
���^r�_f��:�oW�Kdn��S��e��k�܂B�0��JW�)oKR�aA������t<`���״����e]`����R�^�W/u�4�5�������#��2i��3��>�ow�v/d���oX�AH��l���!��E����і�θ�1_n�,o����eڎ�n�Vڈ����Z���7�3ѽ��L���->�՟~��mƎC���En�9��| ���>��m��.��2���21���6��ݼ�L�����Fњ3��������h�3&1H�G,a�,�6.�YZٰD���@>I'3ܳE�V7lF��+�	�7�������v����J}�*�Ґ�x|�|�h��8��s��f5�ST�}9�W&��g�c����������;��.�[*��&�;��?C0Tt?�^��"w-v�0Od#;��#{� ���
�������?z{���8�?툙�+��N�[�1���ˠW���"�H��ݼw���� �v`,��qB���9M�NGy��������n���B~<w�9;�P�ۯ��xi�'�u�aK�Va��������#��aR�>�sآS�抖&N5��k���yydR�nl��,Z��ٮ���8+��T8 ��R��a�����*L������K\3'����G{BE��;�ZXn=�l��w�ނT[k��z0ͧ%��S�Jʴ������v��r�p~;�'��#
�E�0�e���e��]�`����I��1X���.���H'�ݪ���M��q;1��R+�]Qy��^�bN�ߵGU �<bX7'}b��Қ-c�h�*o��j���^�8z��M�5��׬Rk�V�8��Ǜ���Ty]FB|���{�0r!�t��k�$(̳7��N�Q�����<�Wr�x�0�V�]�a��>�}�⬨��[GTi��P�9�
�W0<5���5�jh��H&e�Jc�����<=Tb� �C��y�XV�*��x�jS�y>�Rf�����F�|���l��dS]���'NRv�#0~����CAlLeF�y��܅Sq��B�t�����o1��Jt�H*�v�>��Ll~zeP��A��,�~�G��e�n�r�U�r���VӴm��`�꺡�{Q��� <��(E����1���zڄho��#���-]�xbI��S'�С|���Z9�x����1Ǧ@<���R�
Zr�vJ$pV�D�9 ),n��ǩ��1m°��i���;!�ͪ[��Ov����
�f˙Ah��7>2H*+P������DN�t��yL��'|������j.;y^�2��x�Â�Y��?�9S1���^'�����/>w��"*C�X�7܎)ȺK���8o-�S�2A�Q�W���3Ih~X����7��h��������'�����D#E��$��{�̤��3�m7W��ڶP�y��־o�����~rk��\��Y��}����giizl�ڠ�HZVy��684�`|��v�]=�-+�t֬�j�*��@�#K
�f`R������M�/	����3pbg��H�n�-i��&�L���g2�J�:p4J����OT�N�1O�����k�����|�O-�v��ʋ�m�gi�ǋȻ!Z��I�L	ygi�h�E���JŴ����oķ}a�J�{�*s����^�]hh�c�)um�7�ʕ��弉��s���'V�hi39٦O֋�����[����ӡ�2�Τ��uΛ��N�i�k�t�i	�3�A���D��p��y�谨F�_b���L��7����3z�@ $Xv��S2��DO�+U�e7c�	9ꁭ���>f������u�<C�Pwz5��q��+#LN�hbXXƓ��pSqԲS��缟��z>���f�Ե��	O["��'0�ku�w@;p���;�Uu- �tP�`���.D��.߼+��9�9� <\}�����r�^�޳��f�B���<g�c)gfR�ˎɴ�	at7��;`_���$��kU˼��4`n��[it4)������d.4��z��r�z�!,N�������O��WfM�GP��cE��*��tr���F����o�|��t�F�E�ΐ�2�RFۇ�O�غlMtD�*��J��_',��0�:�y����RѢ���ԁ�]�q� q�
I��EsK�PO`�yΗ `�a�B>gg����yD2(�&dC�lo��d��I>��h���/�#��6���[�������\�1'at3'��]��j�r�D���P���s�!��z��4�%�[`��#MkH� :5@���;�3ܖ�)C��C$e��٦V?���SLQ^�s񱴯����
�xrg:Y�k��{)�c`�E=xl!%O�yEIW��;t��+]RD=��g�����~N����̭_)'���!����_�Fg��L]5��DS����ev��2�!��ܥ��z`�k>]�y���m �hM�|ؘ>&�.��/!ШFH�PHb��u�}��}sT9&�Ь�L�ū'�wT"�'^`a�~,�6A�̔��w�����읃�RM��?h$Z.�_��N��qՙsE�F��71j��qv�d�]��¬@ȥ^�L[B%��b#Xx��ïC�IX����=���������ZQ� >i�v�0�[����C ��?���������u_=��=�vRZA��|�,1��'�3���2���W���2�t�
�D���k�f�l��<$���%bf34	�)!7�9E=�A�F)�~u#��#��A�h�D���Z�a�jF����4#��;�?iB���ChZ����y�ʆ.#7�|p�v��hx���60��Ge�ھ�Ua�n�ǥ�|S�3z[l�0�E��6��5jV��vv�p�6@W�-al,���ڡXH�pu�/���|�B��!q�Rb�LfU�t���V]�{��t�կ��=9e�!{l�۽tj��G����{�I�؝�u	Z�Q�QG�W�>R����� ;�K9MG'S3�W����+2����~�<������p?�{���q` )���>@�t���z��a�_O���0��f7v։�@�K�?�r�a@<!��v����`=�:��;�613aɪY��ҪyԐ���rc�!�O�
�����.��q�s�}�?,&K��������i�+/�x��'�����l/7���p�a\}�	lM�P*9	9�����,�N7g��k_0