XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��R4�4K�=�y�� `�p��k*�;ulC��,�2��[Bm���D�p��7v�H����zu
����w1�V�۰�ڊqݜ�X*��L@)��ki��q���l7�p��=I�>���<N~F�{�N �(�}=?����Ï�G���1$��N��� �����׸W�,��r�cP���(�^���m�o�,F�ȓ)��?����|r��ʖ��m~���m&��FP�C�)|����m1�vm���S�"�@{� �+�
�_�U!m��-�5(���
NQy
^;�!m�7�U����ױ��4�=�_1��тA�|E�����3n�xK��5����6�ĥ���T�(��x�+	�^/����䞪OB�����M.8�0ӱ0�b��A)[�k��9�y=X�I��
�4�������S�eu��u�eG��Ps#}a"'�
�8k�6���/_\騘��x���tg2?U�{�������.p6t�^;�x��o�ݴE-���B��D���j�\5U��V"ekT{�L�i��u��,\��t��o�,����؎����ac B9�9c�j
�o"����^m��C|&���ҕ*m����mє�I�gXlv�cR�*��g��-�$�IAl�<:l��۞�B����_�Shc���gCµ��7spYU����*�D��X��{�e�<~}:�ɾ�G?�a�Or�L�m[&���VZ>2��ii3�V�����ܼ��A�[ ��Q���Be6���7���lXlxVHYEB    17d8     890F���
��cK�Ej�\G��a�O�|:����#ʪ'<��@ƙ\��,��+�װ2L�d��9����s���t;��	o��L]?ц�K22!�-�]}����9W"v̔����o"��y#��n���E��%<������n�揬���-RGF-Nu��Ɇ�e<@$\��㰸���/�:��zu,nq�&�Ӡ�ҖY+>SU݁�nb����H���+(�גC�;�~Oi��0��lg�ڝ�҉��a�W�[�� �'�G�=ë�!��Շ��[s�GIJ���I��'�@���t����W�N0�NK��Z�v��t�}��l�A邕��,� ��X�/b����}��eU�����GOtJ�d[��������|�q��a�6~Yi�+������d5����<V._�G-
�3VC�(�'Mg�S�.S��22t脗8�������$�)�M�X�Z4U�C�e[8�����7pC�,��ڬ�u�?q�T����S��%a��K^2�����0���Â�WG QEa�Xn;�&�֢`��1�r$�	���8��BM#�8v'�G��El8Ô�n���떏8�uJsb.6�(� ܟ��n�~PA>��Z�l/�Wys��3�6�H"�E)!,�j�ܛ��ī��t���E���!�R��u4������Rs�o���jR��U�9W�}���RG���ԋf��=E��K�������ٱ���1��Z��~s�u�����1�\�_̖�Zv�>��3~T�7�7��!%SN�h�d��B��nn��l�(��z��`��;�����!;"�;Z�����'���L3���{���W;���;��fU��+3&�uǶ��bQ=�5"�+G�/���9d`�V���P���{G3�
�1�[�A���D{3��$|B{&�;�=e���ի��M�;��w4�xuG���[M���%��5�r���zhR��b�~��B�������5�lp����gU�ō�'y�S�|i��P{L�T�`�3؝���$!�اrp^<�ل������p�+�`sT?	N ImQ:Ӫ}S��?�2����H��C��Bg�@7$t�?�ߺ��	y\����E�8�9c*e������5i>���_dRe\qyI��y�WqIV�c���L��є���ʝb ['Ig��q>�����}m���D/�ip�5o!7�����gSZ���T��tx�̵*{7��\�3��O������� �ʮ����k[��>|\	}ҡ͓0��]$Kh���gFs��}�2&�>p5�L��q ��%ɔ�t��9E�����P�0�y��fC�#RQ�~V�0���V��iѠ.���P��� h� ��~mћ�/?���`� �9���,
��`O�O.ё.��t�Y����V���֓'7�h6h��(:���=  e��`������WMƻy��Z�^�$�>l�/rRIx#�J��� ���O���5j�
��b���E���W�C�n��{{���C�'����'͂��Z���<��-�@uL:��4+� >�"�k��
�5'n�mQ���C�ٽ�i�;���Ox+݁e����#���n���Bq[Jn��" �n8*�p{�ד��.��@ű󛾑����òw�[WH'�
�8&�=vV�"�s}#�lr^`�
%K!��c}|���ӌvFW�V;˽�I�� �sī�k6\�W�N��je��K3���&
.v� j�D�`-렘����Ô"9����t-�J9�w��N��<��ʜЭ[�ȭ���j���݉�dV>f�'��u�G�2A�U�8{os��y["BS��)�qGC
�X!h�e��A�d��q�����qv�k[�V�3���9��f��>��l�^�w}Tf�N��wJ��e/���ao��?
��*��cB��@#V_�Hy,^'3�(�٦ �O�S���Vr"�E&:�҆N���FO�Y��F�~S^�Tf�2H%Cp1�m#1FӅ�n�9����½�z�6�C����S� ���:��w`fq��U���	N�e�ԭ���͈T�9����8 .z�r$�h�^Ff �
I�:\?��o�nu�jd1�B ��W�:q����U�g������b,Q+=�֫p�e0y�'Bc���Dn<�b�3�=��S�