XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������N3R��"R�Ш��_�v!u*�zoSd�i��#��d��tO�$Q"'�se�;����ٗ�R��#��2b`̨���'�ip�7�ϊ"+�(00��������� ���{���D��S�O�>�ԓ���]^�{�lH�e����K9��p_�f��3�kB�=]p4@B:�p��~��s`(Y�!�GkN��ij�¹�y(�l4V`���bT?;&�G!��s87��|ÿ����\�H~�ZyL*ۭ�Wz*��la���x�3�FUF�r
1r�s�_�S�ȃ ����>�!g6���M�J�P�:��G��6݁a�n��@�;�H�����n�[���PL*_�L��gj����]<��Iz*_lR���h��b�;�����P���'�"�>���W�ʇ+(42dfY%�}�WT4���C4P)"'��Y56� ��N!��w���J�U�"i&�l�^k�o��-��(j"g��0��BE�Ix�T`pç�,�S���J#<�K,�	���I2U���l�[ޫl�͇�/�7������r�S�L��MJ����]�9�E]_?X��O<?�+�����p�}�rJ;��[m�t�^�Xܣ�I����Q�����'z{0A���t�BQ�"ag���-��Z9I�/v%��"���W-a�j���\P��)���1u���>��쀹�b��SMZpl2����]�*Exd�J���c���sz���dnUdl�Eԛ��Ɣ_#�XlxVHYEB    5d54    14e0E�eyc�G���^~f���hE6)9􌗧&��h��A�T4:��bOw����Ԟ����ғ<�;^�����zJ��x�n����?�ՠ����Iv�2a[�우�,`�MS�mN���#�(�ł�{{�]�J�'7@��OE�㳸���K��Zᡋ��	�v�n	�5Q�
�S��r,5��{}}���=�ط���1�e;Y�*7�"������K)n�$�+8�}a�X��f����P�|~bW���  ��X���Ca�T:k�����t�5Z�8CPM7�R�8�<��}iBc���"od2�b�u��Ω�I����r*���&7�e@ǉӤ�k��)O��z�=��2B��ˁ�_k ):5��f�1�g�\%�+���T�T�������կ�'�d�D��������ݑ�Dq=)*���>��*UU��1�I{z>���=��������}���p��h҅�����$%����}�R�*��ʽC^^������&�*tbW�3Q���>�ud	����M
Wʠ�3�,�������lhO�j2�Q�A�s�$hf��Y�E�"4V��n!����z%L�2&����N�|ޔ{��*B���#�B�#P7�Z� ��"�kB�;��[���#P��$�� ��2(ɓ��B7Mz��xrb�H�H#��;�������8���,��:*����0s�F��U*a�a�lէ	1���:�[I���y�:����8�g�?�,�0nZ�.P*�?Εqk����咆���:XsC1���X�AE?_��l��%����^�|L��V�����B�f�-iwI�B�d��a�&ym`os��&�$�,%{�r��n[��������<�2]�"�!�u�=`�Ȅ]��O�g�$_"�!4®b<��S��ܵʾ�ĭ��2�;��+b$(�X�� �Bڙ;x�ٺ��&���I�,��e���]�pb�v�;��y�ɶ��l����p-Us���)3�"��Jb����8�і�|��z�w�� ~Y�63�J̐�4�/|���㺊Z�T@���pu����We'�\��
��P��T����4ɬ�o���q~T<Q���?��O�R9p=��~i�z����������Řn0�}wO@�㉩�IN>��l�I_]ÿ��M�=�/%y0�i�9d�;Evc�;�Q�Ef ��]W��.5�-��ȓ���,�@�3neSI�#��"��^�q�7
�IS�-vy�xZLۻ��߹�m>d>r�%aWK��Wl	�Tm�4?O���l��^+igY��$[���h�c�{u���+�尣.���G)���sod��ҢL�Şk��KV��q1��"��"�e�{.wP�J~��M�!s�X��v&�]���̣km�#��m�dhK�H���_�GM��\s&�߻o�j܎�lH����3"a�u�s�q�&��<Ӭ  6y֢qK���H�C��&:;�i�8]F������}m���-�BU��3߽#S $����Ɲ��UC���g��7����u�)G'�}�t���w�t��?�x+�^�j+�?������D��]��^��<A⬔�a�����H�ݩD)��Eq�F�jXd ���mC�^�o%�p��p"ȆŅ	5ḙ�"�V�B^������>|�<:�����@g��Vۦ�+�E����I|�-9IS���^D�<�rL��л!b��舾��s�{��c�����nS.�ρ���EM��!��q]��>ύ@@� �C;�gì��f�����t��yEJ\53Va�fxu�� c��x��a9�c��x���1�qv�+�>�w��<�qR�<SL>C[r]˹�f�J�v��Mo��O�siIb)L#�nJ�i|�G?�7��}�~Iv
;��3NC��?�"-�a>Q*@���lΞ]�d��SR+*�4L�7~��>���!�0��節Rp�ݸR�bգ*��v���"�w[�:�"шҽ�dl*�w}�EPW*���ï�S%J|c*].�$�3��u��Zu�BF�ZiJ��~b��F
(9em]�s�@��p�<��`�p%��{����8s�1��/h�A��X��ti���̎h����L#�"E�̨�)����%K[���I���T�s�YW��1`6��� �ҋ�r5mL��zT���vpۦ���B����i��ԕcR�Ef5�1Ui��ۜ�9?^{��Hw�\3rҶ+p껎C%A��K,z����)������Ԧ�V�AI�w��d�M���=���5`�al��'�WK�\�pZ$��T��y������"��pő�K$��K�� �� O'1���f�j纒V��s@���)-�)��L��$3��	�b��l��K���(�#*��߶��1��Wf�Mׅ\�?x9���t�"�e������w���~P�K��lg/{�14�}�����.��^0���!7@��Y�Q���V~R���1[+:�(�ůz,�D�͝d�e����ᦞ�V��z���n��Aij�A[=f(�-�R%�K�N��b�́izC^��l���
J�azF�$�^wzD�h:îP�
``�QxQ����~h[��[�W�~�Wj�Y����f��r#�؞�u�Ѷ	\�7p��?�0Z�s*Y�Z�-i��<z1�޻�͟��n�R�h^pZ�������n�!�6�^�߃���}87�\Z+@�����-d	���4/<�!�
���|��d���%$�-ʎ��<㭠�А.�!��ys��r��n��=��yu���	�|�6 +h��b�s����.�OSr��<�9\�ُ�&ƈf	v@ౌ�_Pvym���fGZ���[�����a���eh<�on�5��A�*%�"�#U6�Ij��9����EU�E�)qN�
?��ꢋXK(�`�F�O����s�$�upr�H/�����<���K�q�j�
�=�֌5qbQP5Ǔ�pR~T����!E��[�/�'��Y�.-�C��X�b�|4X/A)�p��ԁ��;�;�Æ\ס.d�sd��p?��\�(�,C�a~��-Ę{�
�A 	E����*��˿պ�`%�84b��B��+�i����Zl�c���Ykė�ɕ�Q���B�"!��-X�~Ɂ���0�V���g>xC�pҥ�-���*	�%/�k�Bٟ�nѮ��*�U��<8��A'�kys�-���l���k����cs�݄�B�6ȉRy�G>���&��q�mw�D��YAE�������TA��u�j>����*w�$hW�hv��E�8�T��^�����>ᄆGF�א�۝�&.7�eI���GyٻA��/�q)���t�mC��/-!b�S������y�.�	!Zݵ$��T�L��ZG�܌~�6�F�5ad+$l���V�j���2fzr�AQ�&�i7�Am����]\��~Z�и��V��ʔ\d!RM@nTT������^Rɗ��6'�̥8�Qv��R�`Q���}��W�;15ޚ��ʘ�;@���@1�c�Ͼ��L��<b��v�iM�4�k)�� 2?8���na�6�;��)_C�e�:i9�0��e��d(]��A8���94�6.K�,�qӉ��ju��T�AO{�(��^�*����Εj50�sC�ʟ�/p0_��/��`T����5�E��E��ηWX�:ϟl�f/7!�0fy�F8���}Ӣ}��a% e�a32>�� �E9%������=g5~g�;"/��,�9��0��R>������J�2c�(2sl乌��U�v���3�m�Ks}������ݦ��7ȩ�K�hۚ
�+�k/{h@�$]��ޠ���򆢀�'�)]jj� �V�Tb�6.Y+���N�~(�!%bp�R��Gg[J Q%�sp��3�[� �E��'�����Q�"tϷ�%���彍���0� ƕ�Z;��v|�"�n��t|��F��
�D-��Z'��9rI�#u��ǔ������r:蒙��9Ñ����@wJ�꒲,d�w��y#��8�(A�n��)H�]}��LbX�-*�t�����e�n����;�C4N�|�>}�~�O5�s�N]5to�! �?D���L�5A���4��? �Tx�5����HX�el�s��i�h�h�|��<a^�P-�nv��'P������K�.q��]0dk�|����$~���
M"UR���L_K��+�`{��Ɓ���� ~�b+[7]oB�T���{s�m� a~�0���]¼4�������|�`�5�`�A��v�Gh��\�P���)FC�!{Nl�BւN���s� ���2(�s�pi{W��>f�34y��6A@_z��Q��=�qRt2�`������<��za��L��~`���g�'V3�y���7?��� =�SJ�Y�]V�|�4�9���Qe~Cޜ��5{̜6~��QS@i E��s�{���4\�ć#R����ղ�-RĿ��z�;�,IguIt|������e�P��|����^�"5�oH��p���-"�NU�8�/�N��`�9O��V��R�E	���	�6|��/C=�:1U�rjfA�u`�$�!L�3jK��)��s'�		,����ݖ����Z�
���z��ޑ�?k��l�
��#hU��͊n?�]5H����X��#��|��ٵ�����i9H9�V`V�pS��~eॏ�b����`pg��W���x��45忭K�TA���\x\�1����),K,Z���זf;�K(e���8���P�suCP�[}
�!_��~�c���4}:p��I�d>m�ޟZ��˼m��RK(�5>l�3-ى��Y�m&�tĪ>�:�����LuF{;���c24E{��t��Y��n�B��U_�el>j��H�6���x��1~� K  �}
M[`1(���� �����l�g����wau�`�3���zy��H?9���u�kh�;��G.����`ϟؼ����l+�������ؾ�t"TVz���rz�qP��^��W����S�S@:C|S�0�Q�1��1� {���OS6͉������&�-P��`�G�o����[[l_��Uy�t�h��Fn~�]0/8(؊����@�zţ�U$�4��&/�S����f x��cx�yZ׃S�wȌ��!<E��)��x\V���ơ�6�]C6!�|����*� u\q���nӗ��-�(����q��Z6	��T�cW7 �h�E��0y+��ӞM�{'@mE�ݟ>}��[|�m��4�tTV��\�A*���|�dL�y���R�f~