XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����m
0�ZF[ˋ�g|[�%+r��j�}=�;��Z�!�}읅��IM���љ�^�7ȖK�w��/Q�D��˯c���kS�� ��	�*y�&��M���ӫ�I˜����8/�i������7���1��O�TL�[3�u~��A��ܷ�g���1ɊJ�Nu��ܪ�=�ʟ<.�y�*2����;�\�ƿW+��K��f�4`HG��"�b��ifak�����j�������	�NH#Y<2���Č�+ދ2zG#�ó8Np.RR4�wʪ��q���ۓ����*��gwUy'�a�e�B�,�tB�%f�j��3|�-Ɇ<~Պ�4���&҃�y��Cǀ�z�l������4R�ʧ4���Ayx�i����
��`�q�<
�j[�����"g��w=9�F�������>̕�Z� ���>����4�sjX}���}�F�K*U�޺�6l%.��3����CY���)O���! 6��,D��S���CJ>�"���M�E��[#���!�r]�#v5�e��"T'3ZDWIͻzY�Ӏ�I���f���L_��S��
ȓ����p���4Y΂왃>��<�<]���߅��k�>��gvY8V�Ĵ�Y(����q�R~�o�O���[����dЯ{s�#�;�N��C�,�s��O�ةܑY���l����!�kP�N�7�0���	�fݢ������{�U��i4���x[$�6Z�d->V�I��zXlxVHYEB    76a7    17c0Y���,^i�r��V��	ػ�E�=�F�C'+��<��~��v���~>羬�f�d�˫����YX�h�rЛ��9�?���������YRc� �nύ� �"���l�'V��-ce�Q{e9f��sE�� ���۞��t ҜQ���=�m��Ύ\n����I���饷Ll4���%����b�t��`���U<���Q�*��Lr�M&��T���2�űg� ����aqz)��T^����}]>�'�8M�k�ʏEx��Dv���h@�s'���N�	�x�wr��Y�ЧV�Xv���k�HQ��f�ŧ7��E����/q:��H����B1�[��%}mh2�J�~DjN0=�a	՟[CI?�s-��h`��;�;W`�N�߆�t�}/l�ejmN%����8%rp�"��Hd� ESE�x9�ۻ��s�a�x�����֏��述r���p��g1C�V�T
F9W���	�Σg���
�_
��8}��?�?�P��J}�т�]�󥓝h��T���)�$Bձ���IF�<_s��δ�C�~�������6b��x�0S�_���Ir�޴���n��2=���
��,��Կ�Q�sw6��H��@�9�p]1>��|��G�a(n�%�8<e��:�/��x�<���洴gej��"�Z.��]]'�t«R^�F���E���_�v�3U�/
�w1�tmeB�R�P�
鰣�qu(�;�nbO����du�d��I�5���=7�2��ó�ԯ,��S�����ԍ�h!"��q�K��%�0���"!�FA����xݕ�X�=�|ζ�g$�n����+@T9-�o'����*b<���p����a�i���P �p��~�r.����+�t=�VG:��7�_���(����A0ڨCG#���}���jl"�+zū���}�J7�@��:A� O"5��6�B(T��~~ras\=먏���C�Kv�����h�$.��{�1@���[�rO6��*(-E�ԉ��.����	����ӯIΑ�޺k����W��C鯙.�D�2��D���mh�VQFc���~���[}����m_Ym���A�;X ��p'ho�㼰�i�\�!�\=�7p~3�/�X�˧���Uo�+����ỏ�$gbw|�XW��u36!�CN�K\K�ĬZ��
D��T[bN�S��z5�X.v�Q߇����Lh���[%�epLPr�<��7�4�aJ>���֣(1�O��X�8�Ff�w�s��o��v�/W�R�KDZ�=�������eX쟖��&p���i��Zj���g%��^{��r��*�2��'Ǔ��ne �U�=:����!�"�8)�����ڸ@O����ۈkD��3*	�����-��G�};8͉�XWa&���Q����������g�:9ዜ��$���������e�� X�|�o{Au�z��Vp�'�a����x��8��D����*�Q g��;;i�D5IN;;a�rԔtQ{������B����7q��N���0��d1i�SG`\�SG�Au��i����)�%�W��LE4����m�TdE%_�*h�p��&�޸�V�G��'�mw�ᩳ���a�Ô��E�Z��sĹ�|`�c��h� ��V�PR����Y��t�E�'zx���[��2�}����iK%�L�h�C@�Z���̥֧���"=����
pn��#�=V��V.��@��DO��9�Kڊ	ą/��4TK_�8���	���eH�f�d��B���@�xA�D������-t�5���62P׎P+���
�6˺3C+L�cw]�O�K4f�G��;Ar�:i���ȝ
��$څ��ėh�6G5���f���յ�N��O^���m�:^/T�B�e�9�g�ȵ�5��t�h��u�ң��(4��H��Dr����~��P`�%?Z���a��ґ�x��}�����?��Ķa��ݝ���������+�K�m�a#~���f���~���y'�j���,�����ݭPMg厨PJ��h8+�W+�e�L���n�)\�O���ߗ ��w�D��=��Y�S
�{%CQ#ͽR���Q��N{�>�f�o\e�r+�:��T�w[6;f�L5o¤�|�8�%d���?�u���W�lCg�)22��2�
��*Q��Z�Ey ��+��r�(�
S.gox� K?¼G��,�Vd��2�*R~~�I�`��,@ �je�0�����qg���x�^�@�wJ��@��P�g=s�.�D�G��4i,|��
ʢ��7�G_l݊��}������C�cl,�%���Z�Ȕ��0h�o�,�+�:X�[�'�]��a^6N�$����柲���]�X�-qu�yr :פ�\[�RnN�(ӛ���͇� �)�S�I����hf'BMy�$���`m�A�d}QЄ��W@��9A6�%vf/a{�^(l]s��\�P���2�+x� ߀�n��D#��7-�Ȋ0HK�]\�T�E�.Ly�H/�l�H�4��j���S�.�|��J@�YY~J4KD��LFG�2'��4�" @�@��p_Oߥ��|�i{��mM�4/�^�m5D�w����i�I�������� �̚���@��/����~�e�)�H)�:����es��a���۽,?�o:�v)R��ǰ�|SȬ��E�%)z����bS�/�^J��mUm��j꣊���@7/Q���#�Q�Z��Z�2Y�m��J�gNg�'�Ɯ5� �Í��f��q`�-Գ��)��v?�*��챭lh`�'����E�6=��lz4$�U��X�ܧl	�d�ϓ�:�]&�4�*�5�#����Ǳ1��S6R����1�9p�!��I��jn�D+D��Y{`�E,0�+d5;J�F6��7��W��U+�CfW�9ͳ�t�BiS�����!�z�"Wx�T��M�R���lz��u	�������V�E-�Y�ӹ�U����)s[���0��iF剛��g��{l&LB:ۜ"��J������&�v���Ѱh�3�_��T$Gם�$�5��LY���6um���qx��ʢK{o�Nf5�ځiȗ%P��V{��ƀ?���K#}﹝X9�\���K�B<Bi�!3M����]��%c���/?��K�dH�RZ�{��lZs��ό�>�N9��\��U�j-�6�l�0�r�NCE��/�;H߰�����|4������\d�uiz�d�ǌ3�*�AMK�7`U�*��KT{c:�5�p����`Q��N�avq������S���!%<;�?�5�4���q������8� ���SHn��Dp�AM�i�۴�*��V���^{P�3��SZ;m�[�]"s��S�>!����;�ֲK��_��&>�;ӐíK+x3sv󑝮�����7��a{�M~�D� ~�
���tC��\����V\d�d�x��ɱ��
�v�}��0�8���©���ڗ�ކ\�e�\��n]�Ӑt���v��ԲM���Q=���٦�~�)��e���jl:�"���7�أ�Wʩ��+�e�@fA�0�3Ե'�����pٮ�U �����!�?�ݩe/�6��==�Ρ�"'�U>��He �5�r��M�	�1t̽�{����r�|�.��I��
E��� ���������V���oxA�`6��	>�e F��&�	��D�HW(m�I�꺗�_$�>�*��
�я��	?=ѻ�����M�<ecd�H��L�A�����%��~;R�e{#��~b8*��j�M*�v�ڪ���֑CZS�y�&z������֘�,���X9��~���?P��~��� ev���W�_(���bk\�*��
Z�6��lmd�8Y��#���Xu�#�)���bq+@-U�����:A��X�E�`�ｫ�T4��,Yl�y2G��=U�4�(<b�ԓk����g}!�ڥ?��4~�)��"1w�k$?��� 	l֒�ɴ\���D�0�h5��.�"��$��mtm���m��E���&�,�����k{ƶq�B��X�1RP��$���N�o�cR�=U�z�Ʃkr���D�BM|ax�Q�r��sփb�@1< ���h�6" ��ۯ\�B�A�^�.�ϱ������PP�C��ʢag7c�<dַ����m��T��D�傺x<��J�͆����!�C+��U����P��aYf#�lP��������!0W���0��`�LB#7=��o��f�L��^���T���(���=���d8��V�-@żI��<�Y�4M&��H�0�� d4�@α���X��H�Y���`*�1u�e}�)�J
�K~^O�M��YW�|�G�����ǡ�m���t| !Z�U|%LE�j3*��[q��;���9�2�.ӣ:�Ֆbw�Ut/+~����1�l��Yz7�6P��
;C���n�/"�����霳���#ǜ�?RGZ��z�+��BD���iX�x�܎ԅ�jC;���s�(�V�R���)x�+���	&9�X� ;4 �]�A?��|$�TS9�fIO������V�xm	�����1���)HPo��KD�.���F���QKی�@��1�����^}Y��E�+ܰ�j��R� B�2����\ �Ĝ�Q	��"��wɎSBއ]����3x�b�{��l"�w����]T#�Zk�Ekv�g���{���z ��l�o����|w^��� [�����9v�a&m��"9=�NO6�gi0^�BRU
rz���l���@u/N��}Z���&��wB+��<����4_b��Im�)��{�Y&ч^h�g$��`�ѭt�~ٲ���X�x)u�A���>����H3so�y��pw/�#j� 00�������a�=�Ue���^��vr)a#QE������Y6y���͸Qi������y�AǏ�gaa��ӌuT�fZ���8{7�k�0DW�V��P3��K�|T������5�Z ���pQ�=���c�f��s.���P]h+�F�z2Bgh�a�o�1ib]H��B[9b��L�nɽ�q�Ɂ�4��)b��*�����h3%:��<c��+BǗ��!�W��p(���B��EN�ځ�#�.d�E�1�l�(K#v/8����A�2�9�	�	E������8��Vx��(�%��S�@3���uIy���}3��cw4�ͶB��z��i�8�aN@�;_�g=��|��dj�j��P�
�n¦�(���j �r�z�@@@���(b�P�n~nki;oq�$>��@�Z	<~�{�y<�/��tu~b(A/�A�!+�>��"�3ј�k�T�ߕ<��]�E��Z���;˧��.]�X��Z���^�}�{�c���X"�Y��դ�>�e8��G����c�ݛcg��t�6�ma� ���z(�5�0R��
'��=��ku��&��'�F6c�۫@���`��Ģ�0���GI�P�m������)�}	Bb/��J#��G��E�Lj
,lE��?a�d�͡X����5���o2!q��t��t�
P���ϔZcЉL	�x�oE3�}��HB�jEW����^�E�=��q�{��d�v��o�w���0�W$��.&z�o��gT�0}e��G�JrSq��ȶ���������p��G����E�	��y��-��y���L�j@��vy�B�'�-5áf��6����W�.&�����rؘ[��Μ��T�	�,��� Jq&�7`$a��T\�>%���뵓v፤��p�I�1X�r�BFuk�7��Ȫ	�xTQ7����VG��|K�j��|mF��K^ |=��-)�ـ;H{�C7�v��U�^�>�i�ua���/3T���J�o�^�0�)h�9���n��'R>��,�����nP�#�|��أ��[�RH¼d�n�8�c!�M�LJ�F�)=�돋p�.�*�\����P (������-W��K"���� �'oPy~�e��3�H��