XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������҅���~8=����$7����x.��>��1e��F3�Kl��^h�:8��]\����3]�!5 �fk�4�U�atoT�Q�k��xp��{�����Մ���gLd\i�J�Q����=lU�s �Y�ts�h�y-gp$.z�C�>�����dzߒS�����g��-���x��r��n҃�Bm���B��zJ.�⯘�?�����
��tg>��+|N���o�N��0ȕ���3�^�4}�2�Kùm�7Re/E�Б98���\.�?� }¢�0��V��y��l[��cX��~y�M�"6�Hv̢.��v���4�Y��Ii@�������/����U��q!��f�ud��.k|Z��B�G���
������-9��:�	��ܫ �Oޝ�Y��T΂w.���K:~�}lf��C R��ẃ��®�2��I��o�b���]J���lF�;��`�����L1-�Eh�=s�@`}!_
O��Q֘���.��ϰ��@�Q����ރqٴ;�·��?� ©�[�݆Ih�:�#-f�*A�JT� kP�D#�t8����(O�ʲ������۱Yv���YMi�m��}S��Xe}��,=UF��iD�B�7vҰ�Cw�A\��U%{���']��F�:U�S��-3w��1!/��8�A�C���l��$����H"suKPg4��Ӕ8*n0
�O2�� `x�Ǝ�&�)?|��J�A˿��dy�0���>4����x:'�b|%)�� bXlxVHYEB    da59    2e30:���d��<v}>��F�Ba!ؚ�{0K������@f���OB��8�_D8��$[3ڤ>=G/�������BZ�x�'g_�,�u�n=(X���=�z�,Ύʢ��8���y���k�>�4M��}�����Ʒ�}� A��K�� _�h rX��� \��-1	c.�����M)Q��f��� ��C�!+�`�Tz����|�j�W�5��,�+���x[и��K���-�����q� ���j7=���	b�}L�Yl�MW�.5fHX��}��E_�R����fS���vڊ|�)�6��;��}�sn��9]löO�Q'�J!��r�e�T����p��"☦��}SER図�6).�[x�E������7�jG;�
p�_�fd�2e���wq��P��O���i�U�1�q$�`�9�@�sS����n#�&�`Gh�8f<2jZ5�s!\����W ��w�꺱�La�����+eE�i�![Cs���J۰<���(��c�9)ؾ}��D}):�0���pj)0�)��,6]&1c�1*�!ޘ�6@�� ��E��Hu�O<��f�`��r�Oa{Cv~�Zj͐Y[-W���mJ�"�P>������<�8��]@a�i�F˝^�Z�{��OI?D�L�_ʘ"��^T�S��e)o�=�@Sb˔0^���S�8�ʭ=��g�<�����Ιvs[���������� =��%�j���>�Ed�#���-�5f��R�#$�$�,������pC����m��z�5G�*F��^��>@9�o�(qۻ��c���9H.��Q�' N�9��E��9f���dĘ\q���GM��CW
�ڵ0��qO��z��T�6�~�~�&P��i&j6H�ș����'�3���iLׅCG���PGQ.�|��C��,x�[hp�\VJ0�G��)���9	[�@3e�Dg.>�w ,LMSrK���s���5��c�н?����W�vU��L�G��'e��c��D��e�8�g K�x k�6�Pq3x�bM����3^��=���2���=��I3h2�븩a��a^s*3���q�I�#�-4��1E	3e3A�9�S>����&��"������3�6T�ю˝�%=�J =ZM�/�ѳH|��vX�W��U���%��z��M�Z6��z���C��ߙ!�R�uX��, �]_�h�xM����7��DC�V�;,'YN�����JJ	� �?wm߹�Ӯ�Pt���%�ԥ�����ߠ�!U��[�>���������E��啧��Y/�c��廈5#�j�F�}��kԪ�0<���!�������mQ���gY�֚2�H��q��Ȗ�K{��a��r�W6�2c$sh[c?���?}�K;�vz��?�(��k|UZ<x�(hH��o�Nm�ZJ���	2nR��Z���HUC���Ye�<�C]	��:�� ;<���2��d�Y����$C� l��G.,��Uu��c��~;�����B	K&����4v$:��i�P𻭄u8X��A ��Q��������(��P�6����ZmKVZ
52?u�Q�l9�ӤP�oI�;m��${�{6����XSg�\��\p�����ن ��`�
�@�BeҖy�	4?ͦx��B�z��=n���pY�eO���������3��q���m�\T��ɼ����w��0%";���+�7#�����W�	�N�P\e�iGᓼ�?적��Z��L��Rl,��뾒�wQ�B$�9\L�㮒_ ������.Y7����)�?W�E����+���2��1�����,q��������L�{�׿����Z�����1�-ʧ˔S��F��!5�oW}��G�S-�ss�uAAi{)�Q��A��	rуR�����)��	���b�3~=��#g�z6,'�F�&�_�i9�^��.[�z_�M�1q�[j�mz�mU���S���J����S��=~��ŷ$�WA�D��y���nFM2�R�k�����"�VDt td��Aۡ��5x�J�!?9S�c�k����7>�,P�-N�(��`N��?i{"W�]��ׂ�}��a���o�<=�}^�q%R:
���K9����|ǘT�|�z}�`ST�i���r�x��)3�Oc�p�5M˂���\w���ٸ�5���1s�:��W�`�C�}�����a��{R.�I��h��8�Y`x�F�@�$6�S	�#"R*N�G��է�lc�m�Yq�袭���Ub��P=5��b1���f�_����

,�b�ZkΊ�+	��'��v0��J�L�AeRT���l��l �!�������T�s�a��_#������ ��KX�;��c�3P�������i)a�8�Y�x�w~.�9j�"�+{Zj'���F�O�W�QٖWv�(0O]�� �x����}!���5�'vd��9d�����y5|_w�yۛ��tQfM�Q؀�<�[|�j���:��4h�zIN��Db � &߸l�)�et��-h�+�Gx�H�w0�g�u���� � �����o�K|�+N�z��V�6Uk�C����r�LԽ�W��Ԝ68f���xn����S�Vם[�KE]2���Ywd��
��IgΙ-7i�L0�{����vsK�=�5����p�3�:Ȑ�ײU��Wc:/�VV�=���G2�m��ϕ��;���c0�I�闻�]��kW�2T��q�����ٓd��k��Շ[2��6_���@@ /ҫ�7^�
�`5xH���������E�/%�E�b�B`d�Rz(�pJxe�#D@f�{	�s���=&���?����.�q�d��5j��D�Ǟ��5 �<��%l��4�H�S��5c/d�t���MSnb}o�hKA�;*6�A5= ���}@x.��"�+sIN���?��jnHY�H�<�P�z��8�?�`-E��W��6��``�]NB�9�oC��v�"��;�c����}������R����A��[@�hlK���<�H��?�hV���er�9b6�=��?b���>Z�O)�m��{#�,�3��u���*��&*ĭ���Wj���3���g��e�O%��+SuN��[)��ӝ3C���� @�N��n�(d�5�_K���+�-��*�9�#frްy�Hg�൝��H>K��>���,�A��MM[l
7%>��w�۸Ӆq�<N��Gl@8��D���.W5+;�xB.��ӆ鶗�n�Elv7�a�+,��c�h�[����o��t]T;;���c]F�ŋnb��F���>w�A�o!��,�O�z!�̝��4�C$9�U3=<�{]}>z9����S]�:���\t/��.������� ?��ȅrw���ڛ�Im��+�O����?&aR�ä1�b8(�i���h�e+���+��z��>�%��`Q�[;cӱ�xV/���-�t����`oف:�	��R���ޤE�ε5]r�.���xDN�cEWj����R�%��;��0�G�B���t��J�����X�Y>�>�?�W ��l�8w=B+����C�ĕk=�k�4��:��8���?����y����^ϔCa'y7���${�R&�� �ጶ�L����w/�u���j�ɑ����쉟C ּ�R�F,�ƋӅ�����ŁP�Dm폓o�6�Qw#4�A���'	Lc5&�"�!�Nύ�N���G;��N�m�)(�X]y�º��D�FuK6�]Y���2�:�SH���^�I�yZ;���L� �� ��b��=IJJ< Y\X���9:@�}&_�k�p>����5aHL�ZF�}�H,�B�v��V�Sw�m\K�:oEh�b�_��.Г�{�]ea�Y=��?n+"�x�N�O��Pn[,L��Q��-í5���>4R�_����6��*�n�V� G�r%)'�H�b^�b��ҷk��0v٘�l�����脶��$�|$�����x�@$܁��2T��.��{� x�Aٜ�����1�E�����V��D�2�샩iB9%��?r�A�δvY��3�Tw�,���K v��
L�����?c�U{9�`�"�݌��\�ʘ��#Λ��y>�t�bF�W̏�(�(����m�����0�1X��%�ߺl�4������ns:�}߸B=@���t�mc�nL(�W�e�g�_xP�����O����N����"'�C���`$k��5n.$�S>goY��sKO�Ԇ�j��9gD�=.)\Dāځ`��K�C�`G�nVm:��}��h�5�߃���l���9<�!��?r�kA��W_�����8��Q`S#&k�=)d�tNY:�8�-�l���ԙk�_b;�v�̺�T��l�~&xL�Quz��'i�ݳ�zwZo)���o��"��M�:'w$.=kx�||����@����j�> %ߙju�u�f��G�:�����u��R{�sA�['{g��ǣ	�j�M�*j�"�|��/܀?�������;!��UL�%����Eo��(�[�N���W��6�XR��ߠ����|߷*�M������f�t^��Cq�:���(�9MC�k=A����W}�udZ����]T�r�!��幧EA��+�S����(����4��b��yn �M�:VK���{�D[��KpE萅��p�;!�l�lɅ�^��\�
�_Ė��1����>^l6������/�κ�YNW�1��O-�E���X�X?f�a�O;/��n�P��T9�:�M�����Я��'���O @ >��X�vM�R�dA�ֹw�_֗�w�Uǳ��rv���A��zH�A��H_T/�����Y����lJ�&�Tk;?Ƕ� ��i�0|G���\���f���� 
7�c�����Һ�Y뚰/����It�$$O�'Å31�����j`�hdq�tx�b�;��I�X�I�70���M�*�H��ef�.�gۆp�3�LE!# ����\�Mε��;J�!b�̮���u�|��:I�Őm��T޶n��	��7�RO�?�7���>�u�c�kq��ה�j��Q��:@�P��A��˸^���ݍM�X`�����7���=�w�u~W����{[�v7`&/�����(�qw�_y�+t���/�9�P��)��e�D>�QZ���@����THg�/�.�11!V	�V��梹��P�ߙ<����5�mğ#:�JP��B���U�ѐ'g.y�t"*A�@g�ΚT�ۦԶ��A�Q�����s��*WI�����﹊l6Vu<��N!��l��#Hn������v����l�w�G����Rx����t��5_v�Ru�I^�J�ԛ�)R��,#J�r���(Y*�/Ҙ�֙7��v�>o���lU���^�m�h�xN\z+�:.��2Z䓛Q�~��ި#9�����i�)��Xm]�qk�*[�)g�{�mN~���0�-��܋y2c������=�1"�p���G?� j�����QhU�	?I�y�	��F�\ Ɯ/�"��W˅��{��=�ޣq�X�� �0�f��y��l0�_[�Ȗ�+�uk�8c��x���3���A�@�@5`:5'��9��T�@Ӥ=�X�ʍ���98�Z�;e}O��1i��ʏ>��}/ޔ� ����/l�#zo���:d纲)@����\Mh�� �u�F(��z?�õ��k�Lu��{��=Seq�w��i�=T��3z�6�pWm%�#Q����I�,%�S���e�dVyB�w��{-	��J ˸e��1)���Rf�x�UmyQC�~�Sx�/�y��=
l:�f�m��� AA=<���Al�xZ�kM\J$�T�=�})�٫G'dnS�N3Y'�r��k��y�D�
u�B����{����"%���8��Qk�l��i������,�ځ����q�?pO�;R"����İ�;T�b�di_"
 <~����t�|z"��$3{&U誩H�<�O�+	QZ7eI���HfTr� ��l����n0��?FҌ�-���?�_S��6���9�13'��EN ��P�d'��`?�y�Vi�J<�7��`����)*j�Z�i�� ��P�q�5lcG���JO,�$-H_���V0��!\��o��W��� ��Rkv%w�"5�I�:=ՄYza��=b��h/�G��^���#� Rq@���� \��P��3�8Z,�o*�;�i�1�\���f��o�D�rk;~C�����i�D*A��b^�X=�vLEY�J�w������������R�$���t�ֿ��r���uMP�^�`�@5��'��LO�K��g��*���2Zgc��ũ���tB�[��h�R�^����䛙e�.v�v���N|[U��l%dR�E,Y����&��������Q���ϖj?���Dn	_H�J��/feL��q����5t���d�����L�����w��'�ᰟ/}�y�"b�j2�	�q��2��aX��z�2�XTb���
X�i�?I��Z�d:=�	dS��Wt8��<�׈�|��B#Q�y��9�(��.���5Y���	Mȣ�lU%���Y��ʥ9�S���is�{4���u�v�<u9��Iw��{��Tw��F�\噯շ�V��w��W(�Y��,��;:����)�H�q������Qe��@��<�"=Q$N@\o~V��
�6O�8����Edh5����tf7����!��&7���_7�uDP��s,1�YF;��~�����HwT�����Ie�n��<�`z�w2�u��<����M��#,�0S�� J
fBF���Nm��.Gb�����6߃������2�޿/|M�<���طX����ի/^���oV�Mb��R��R�0nɭ�XlT�/Q����*�/jU[*�K�	��>V	Ǆ�",����ow�-:�C]�e�'0�� P� ��r��p�	Ů��6
���U���[�i�8�nmUtQ��uTb��V�5>Q��69k�䵀 L*Q�lI�-�'���`�'#b[8�@`�)1������{u�z�Vߔ���?0���������a��L���� �@�r��!9d�z��*NA󎞚�P=>�ur���3GkKA�ܝ�֮ݘ䣂L�θ�F2��u��W��Oy�~vs\�N
*a<�h��q'�aT��cn�E"N�+Y�(����4U��載i6�6�o�Ȯ]��?1���2/�gg����[sM����D��)?����m�܎R��t	���e��]�����\���2�r^�"��:Po_]�M��'(�`�B`O�o.�v�
�*�2^'p�l2�G�[�}�������.Uku��y��m]����R6@{d��=M�=~��|��ϞYK�,�|X���Q75�w�&�����^迨�"
� #��Y��Z�Xq3rp�V����o��Gb\ ���n��/��2Z���
 #��M������{������H)�'�i;��<QLt��벰P�%'l�f�3�d7_٬|���m��S��	���dP�}<���yu'j�Jx�CjE~PyZ�eV���'P��?r���\,Fɫ{<��1�3t��q����S_ �u���[(��>���-�b{��f'���9��F�X/�#[�:�d7�ˌs�:�I6Ԯk���ߩ�9��y��m8>�g�[ؕI�q1�`��Y��i���<x�]�U.#�;�[ �^m5]t2��#�_Y���Rφ�f��mW\�9Guǟ���ط�[��܀�g7�[�T�V��{ڟ��[~�2�~u��	C�r��*���^�C��b8�)2,��U&|qZ�	C�*�3��㶻��������?TZ�ƛM\�辳�W�����͒l|9�A�$��tп9@C��Si�nA�4,3�i-|v9�Y��SnuCbU�>�YHyKV���F$�lS�" (m�G�_�n,�=q�J�|&T�Q
K!^^�"(T0�Ĵ\�1 )���J��"�GY�A0 T��+���N3C勳:�K��vCҧ/c�X�u7X�3_a�Z ���_����&e���gX�@�����t���m-?��ՎV��/�"<k�Z|n�_�"��姜�c�8��M_��5*���� �R�X�{l��@H�i��K�)�G|QwI�m�2����X�7'�V�Ѩ��
2�3D�� �����<�}Q����m˶XՕ^�h}-b�q���[�|ʪ|�_�dv褟�=�
X�G��+��ggcE֬w2������(�	(
J��q��b��x[~����	�kbW׉_�/�Ȭ� Ki|D��t�c]����`'�b���_����J;�#��L���nϲo�m��� �� F�ݸU���-��Ŝ~ʻ��O�q�Y�\���;�S-�����F 󹮫2M�j�r���^ȩ��g4�{����Rj䂏X�V�״e����<�PZ#7Y�D�
�b���闾LQ�y��2p�=s+�`|/���F��ޜ�S�t�C^|�L�m��,vs��Ջ�T�a9��Ipd:�f���Sw��� 
]_J�t�l�f��U-���f�(�F�W��6:����'ǯ�K@�q��(�+��o ���L���`	9�4����js�n4��g]S��1e�W����/����Y��&�(0W-����޴�Z���e�H���$2NL\���P��H�+R�!��R�f�5����z�H�"��'��V������>�>�1~������Cg4��₭λ���~�^���P���w
�s��a#gv	�rԲ��������c3J�F��G�pw���H钍�胊��&�0��JA��H`NE/3����ɴ�"��T����Z���t�s
���8�a�EZ* �����)��N���G���GRj��ց����� �v�R��#����1�S�[��4=�>�	��>�4��Z��E�vnr|%�8��(�7݀��� �&�n������z�rX~7]�E��y���&L�ڀR�O��`9��P,����}�j�[%�~ɨsA�j�R+}b	�lDOm���"-(e��[a�hg��,I�8������Tб{������h�M�-܋� ��o�dHmPY"nN����?��,4�R�\}߸�����WW��<�]�&�$�fF�)YU��,:��t4^ۯX!+t�!�)z�Y�}��cy< ����*4D#�׀��G�F�y��ػ��5&���E6�	!�p ����H�$>��@&h�k���4I3�0���>���בh��Ʀu\���>͟���=Ȇb�߿Ţ���7- ݶ��`���&���k�%Mێ�V���ʬ�]t�_3� ����Ew/��K�2�8ɶ��M�gr0�IҜ�UH/U���'5?�j;j6:�?RX�Ͷ."�,2��	�'�rڿX�О�,�� �CD�c�/Ð��F�	��T�Y66�)��!�T�4� J	Y�Fe�o�%N�#�ۚ֕�/�]%+�`�����"�������r|9<ą�޺+��-���Y�]I}��abS�+�­��n[��Ѩ�T�cB<���	՟-�^��)����C�Q~�l!��g�������A��U�k[[�pS�x�3����� �V.Ad�vZ�o1X��YC[�+�z�H��e�Ή���̇���OA�q]:HZ(r����!Wp�u j�����l,�������R��!}ݧ�W�MY���a� ޝ����7`�A���J�?|��V9��C|�\h?������w$&�����5�4]���.w�%��}:&,�MD{���hS���f��V���`r�C�ӹ9�K������t�=~���~��y�&��	�D'M��C��˺J�n/q1PktF�C�� �*���*�$�;�z@|�!BAs��]{��/w�伞Z�g�xի����L�3����}eҼ�6Uv��`xHK"*b�rje�}�����'yp��d/���`�R����{�R���)���q�f���"�r�obG����7��[�+�	��G���F	q�o��d��%w�@�}
V�N5�,x��,�#^��܇9���r�[�j����8��������q���j�E�ڴ�vx,�&m-�a��/�� �m���9�"C@���� ������|a��hi�4]�4n���6ۈ�k}R:1T�7�Lm�P�@��._��5ٷc�d5��o�ph��Ot���W��y�W�+���1E��v�-�}6�V%"���+v�@�!���hg�$t)���OZ��P�nb���fH��Sw>��a���$0ΩAs���h�L �E�PB�r���m>|H�,�?��A��'�:�
Μz�iUv��ڭ*���aу����X���]v���눶t|� $�Yj�n�B��P�ӽZw�挲%�S 8���k�4&ɉ(��K���5���v��R��4H�1�@zH�
1gy���� ����M��hY{R=^���f�\E�˹밹12?n���ՎXކͪʈ	��)��''9��I�Ϫw&�x����t���JCi��� Eѡ��W�%c�55��0�ŲY�a�2d�ľ�o��Lց8:CmULpz,�;,��<ŲF�P��j`0�߷R_͕$��LN�pC�G�����؇�2���ML,䒫�2M��e�)=W��.4$�;�7�Pn������Ai[����̢Z�&A⇑���)��^��u��CX�ɗ����½kp&vXt�]�,�ޱh[��h?�	Q��0�B�����^
���FyI�*1u���|��b�3{=��]]L�� ��>B��t�L�Y��Rē�C�=��Zn������xd���I��a�W[����(��Wb���A��Jx7�O~�-
��r,�/�?8�3��c��\�Eh�'{i����dZ��%�ڭ����
��^L�p�/ʾ��#w}]��!x��
%	~�q=�#�A���6�a���@}�����7�4�Љ�п�4��[u�2�}�L΋�h�Ԏ&9�kC�(ݒjU��w<E�b�Z<��MV��T��Q���� �)�1�{���H 1��\4���l�c�6��n�|NHH�6��u��0�,W8���*O���r�rGb�G&�L0�'���A�ESZ�*Z�myT�����F��qr��i��i|��pt��U��֊8e�g�L8Y_=A��Ju��XX9�	��XdF
@N�}���e���*7�ͮ�KAĠ鏺����0e��%"�p����$M^��Z�l� �pS.l�*��eb�{�nEF�� j���r�\*3��I_U��
���;n��
�./�j��M�ZKU�Ak���Z�@�0"��vK��Eg�ܷhm��W=G���zpT���ThƤq�����q�JݏbrzD��5�A���I��Ojw���O�Al~�IF�e������3^��<�!�\�[��׃��h�J�3���n�OLl"����z��B3������a4]�o�ەs�GNfC�_m򃲦�b�O��B�l���z���	֘a���Ix^�͗|�3�����Emzb��N�5�V��%�f�yzj^>���K�B����c�^��>g��@ռܐ���q�ޗ}a{Yr���3��w!D}�̩��R�ל��� ��ݨR]^��H�C��