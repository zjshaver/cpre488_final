XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��gX���SN�J��"A@<��	��DC!�m�b?-��EM�`�Y
&l
�G����Ur����P-�`�z6\��mrk�̈́_��S^�n��W5U�a���pGtI��#{� ��Z�?�.�;��F]
�<��H��"�ˤĮ�xI��xQM�>[�b���s��A;9�>�ׅ�ߤ���٬����{6�ĆYau����isH���8��LZkWASE���d��h^�<Q_t��G[UM�_A�Y+7�/��S�m7_���ɏ���\��Gj:�|�K�������X�N��-~R���⠫���(�P&�5��z<�����w4���;��A.BW�}0v�IS��M���*w��8\1��z��s�p� �ր�6j駵�N�X�~;��{��⸹y�z�F+6l�ó 0�Lˬp,��h]za�ؓ}&y��e�M��A�袹\-��ɵꅇ�?1o�}#T�o�;�p?PKzFX A{�de� C�F🫭�R����|�� �3a�i�3�w���Q�>9j��C�#2�8�9�2b��P��,Wum� :��r�#�'B5���4$D��z�I���P� �y�Ve�
��=��f�sY{��RP���-4�i-؛_.p��Ԡr6�P+�����	���?�q�E4�ʯ� ��UKJk~�>X�@�O~P��� j�����W)W�6s�����V��dl�Ċ�?�=�*��OMW�3S/�W�-���O<Y��c3F�Q�@i��P2�A�`�z�&�XlxVHYEB    3da6     fb0��m�X[��WiKn^�n{H���8��ޭ�D(à�{�Ԣ�#��|��O8(����dS8])��(�Л)N��XT�]���VE�` :>#wϘ�QA����E��p�����U�ΎX�����I�~s�񥯱���0��ɛ�M:6�߻�v�v�Q��:}&��x�*�^?7-���E�\T���XJ��e5Ұ�I��}/d��}����Fz�	
�(@ �`7(�w3v�̭H-��y��dC5�'��2�LL��y��N~\"�#��Y��k�e��Wg�r�&��nB'��t���~2��5��<d�6��n*�G��I��� ֦�Z	��	C�N441/8R�%���>ۗ�S�f=Y�� n=alzM�s!��`9�ь�#�נ����q�p��u�
`�ޛ$���D?� fZ�)1�{��'p9�iǞC��mCl1��* $�G�aF�2�`Z���^�"x&EV՚���{>�DuDG������)����������ړ��-nd��x�>���oO�#2|�X'u��ߜ��Yg���\�K[�'��8�_�<�.�`��S��~Uy���d&v/�w�lǤ��BVD�� �����(���=���~S6^� 	δ�g�Q�Y^^��<�)�P����������������}��q�]�r�	��󀋰Ů|�.wz=����'5L�~]7�5�Vj�|m@_����#F<;�'�b�zn�70������lXSCp�8-N�S���I��B3�\�	�����yW7�v=B�ԶX��9� ��4@�\�ߗ�̻�E��a,9�
�P�4Ӱ݊ͫ�`�������0��!qe����:��]Zݣ������AP\%��Lv��8_���胏��?�Sm�:�>��F��?*� \��**��<�y	+�<�H�߇9 �Cbp�
]z� ��
ST�Dа��/�t�x��j���,���^/���|h?�="bG8Bc�u��9#�4�Tȗ�zN�$�1{�0T�9r��R7()uS�B��V�� Y��t�{�J���Z�d�HV�	-�u�T����U|��u�F�
��9*~�i��Ȏr�6`w^e�'����Bެ��F���3'1�U�D!�P{���x���<ze}*�5Pfx��y���;���{c�&�����C��g��o�P\�a!�Q�h@���o M�\������}�ގ �<�5:�E�XL���75O����k»��a��+[,��^ˮ|wh����ʦ���N���z�
{�
1�\��+s���2��ǘd��Z�[ά����0�_�OU��N%���qG[��_�~\i�R�z﷡	��i��_�Ipm8��F������q�v��x������5�Z���t	�b��%PIc�����5Ç	9��"��V�K��e���,w��4�H	aM�E䵜��'B�#��N���5y���O��j����%��lA��������k�D��޵eyV!�s��G�����m	�
rg5�]�������&��gl�����gP�R�]��we���C��H}J�hj����WqAiʏ�v� ����f�l�筌��E)+ۙ r���mS�J�9��'�����9	��Vj�Ӯ�C ċ �J,qG��XαS< �K��K$�bU���E�,\�ߐ���c�f 7�@�x�?���DIʌe^V�d;~g7M��\xF�͕�&�O�fH��Q4��v ����:��uޖsΡ2� �~�0�yl���L-��ƘL��q���E�}��q�D�#8ۨ�M��,|D�AL��X����$�P�<��-����ċ��D�����JN��!V�)j,98�$�]E������'
a�=�����Z
ǳ�.U='s����� j�br�̵ ���&ۀ8�]���n�A�L�4H��oa���e���;n��㐅���"N22�z�֓�r{Y�k�03ҐYn֌�������R
�A�/b+�.� k�M�G��[B�𸇸��:���Dm������(�8���������\|2�GPi��Qf���a��?j�'�� ؂���HaJ��&�3=�ߕ���)һ��
A[�8��h�R�4CUiڶ{i3�S$r��;��Df˫+�cq����yɆJ����in���QⓋ<�x�R�o��=�u����]�Ӗ�����p�4?�0K��>[��e���\��Y� 蹸�:_����tԆ���Εo�*�@����X��ΓVm����d-�a	��5��c���H��/���\(�pm���erX��z7��|� ��1�U����w���|1DC��%��!M�F��� b�D���bJ�KF����ϑ�1�X,M5K6��rS>M����jL*d�9���:��[������ؖ7�:��J����(��J�����"Tښ-L�+�#�]�uR�c�=;\���M���#��{EG �)��E.CX.�|�/!<K�T���{�3����������c�"���V�\P8~�v;�5
%PxwX
,_a�(��W�L{��]�ao:$0m5�=�����֥��o��4�"P�����l�I�.#Ϊ�DC�ԝ��쑗m+yKf��/���G*��ٹhS:j��G硰���(�a�Ⴗ�A�^$�V�kWg�&��G�	�:}�,s��)��r����[	#&��d�,e���L�}ǜ�'4;��R(xշ!q��5�3��G��`Ś �4]� eFz���ɜ��	t\X�l< [3� %$���_��FH��VW��i�'L��W�b|�~}�Oy��F�:Fލ��|f΢j���RȀ�W�p�C?۷aC�Q��v��֝i�x#��س8�&������?S�������˷�m��0q�i���Ԝ���d����,+<д��U\������
��p���4�e�p5���#kI�32/h�����"	\X��T� �]��w���ym8���u��yRDtd����۰���c���h������q	�o)�>�u�F �������6�/�i2�Nhts��>$��F�4�cO��=���Cix��ݲ�:��(gb�J[�ӏ%P�\Zv�ꇓw�]�C/�,.ւ��.����s~ʬa�T��Ūf��?�X#}'��"�hY�{����=Z�(��ꔏM��UH8=�Q��	{��bJ`}�,� ���0{3U���"�h"�H���$�/�G��`��H��51�ɤ��XMbs?�$��͙P�J56�p0J�?�!I�@s=#���nM��:�r����r$��:�yz�M"JR�t�d:��6��(>�N�=�&K�f��T��7�F�1�Ib�)�C��qI�{�V^�͜Ȥ�������ڠKz:?6�� ��V�����ɂC3�:���`����<��1E��EJZ.��2 @ۡz� �	���_Tx�Mm��H;��4ԈB[f[CR����$�q9~�z-�f2kƏ�b0�,PFA���(v�H��o��o�%����<����.����o��-����oh�}�����q���ћ��a�E*�]Nr�2>����u�w�ű�v�T2�.m�_�S�sj��J���w�1N9�Jt�����R ���5m��E��˿� �4@���_)���!6@��fU�$��3���M���me�����5r�7k����r_XE�j,��	LտA�m�N�k�����c�_���J�P/�+�1��,B�0��p�H�7�/ax�R�	�P��@~�7�َ�ذ7�$�!h�`�|\���T6;����:t�D8�)n�L,��L�q�Ϟdm?��I'G�O�"r�">��A���-2	��Bz�^+�	�@�T;�_,�����@�6��n��5w��ꠇ��?<MJH{��¶f���d��U�����H.���Sq��D@,�[�'����Yg�uެ����