XlxV64EB    4283    1110TB�r����:�����c�J����,b:.���9��q���N�����HՅ��p#�T/���*��j��鳳�8��ab��x������M{)��� Gf�2��^�o
;04����b|��Ӂ�읪0A��ܞ�v�_2���|r1���ow{�*��gs��������V;��l���Q��(c_v��jޣP��_0�]�Xq�j�4�X����K~�5�j��F�E�2LD��Ə������f�I�ܓ5fozS���Z����8d��HY��g=�uh7H��F��]z�oJ���s�ܔ{�΅���؇�F����R'@����Tvs�N��hg�<�➣�̦mكy�J(�C
��0�P���@�C�>nW�[��SRg�^��/�n!��D%�O���w��Z���Q�^&{[��.�g5 2*�5HW%a~bbki�B���������Y���)��PAY!��yeo��F���;+g��P�G�/}4��L��J� 3��C���r���D1�)o��W�'�6�:��P�����q�x�^Ǖi��:ϵ�ήk��1��3aRǎ�e4�Ihsy�	p�X��PTz	�H!0�9B�P	C�"y��d�g/��!s�z�Z3T=|nx����L)��Q��c��ࢲ���,>�[�?��5��ȵ��z ��l�ne�؊L�����cF��`�	=S�{26 �s\�E�rFB��Y����2D_�%�[�'5��NRc]��v��J��Q#;c˺� Q.�	�)��*kl"�d�j�kE3M��>/����NW��������z���z��b~�p�r��"��f���'A]�6(y���R�٧h���2O�a5)���T���I [ �т-g�CV��nN?����2�`d�%L��<��[�b��yb|+��F���+�8������{������'���;ʵ{�&���LH�qYxn�MV5|�P���`�"g%�TA*)�ΐ�Qy��8`�!4 &��yP��?��wH���h���t�gM��<5�<�dr��ݺT���e^^4�[
�S_ީl�'W�O#0+���~2�z�Ě��x�AV�T���U����p�$pQ$��Koi�$�>܅�%3�3�.��P��w�/S;�k	�Y������3�8��
�{]�����m��J"�ޝy����K��l�w���SYPqU_H���XA�u_fc;��Uʒ�Z���K���R�-h�Q5٫|��0`�n�(f� �IX��q/���|��vc��ɰ��.6��`=���3The��N�ɳ���{�(�N&��+?^H�Y'Ae���۲w���F��#�(#r"1[#�be���	'�b�ϷNet)O`��ˬ���\�#�p1с83hv�sN�(�c�rG	g�!�9�	��u3P�7����)Һ��m�1�����̂�����b[=Z�v|�Y��};���9��-��`bL�*U7�-�����'I'���"GPOU�_�F̀Z��_E�d}0�إ

�uP�����Ib���A#������4��g;������`4�`ie,A���k.��0���7s꠺��)��M}w�u���/�cXޓ<	��W�g���+L"ֽ!�F`�e��?�?��=2L?$��'+����j��,!��Mw8N=Ǥ���ȷ�*��:o5Cr}��n�%�c��`���`�d����Ȁ�7���k�77��~T�t�CJ��f���TV=���R��CՕ�2ၯf���BQƪ��詞:MWR��榕' mG�,�d2zfj���`x���3i��~��4�?��9C�ֿ0�z����h
��|
����Ќ㛷�AG6)=ql���%>��������j�na{��64~���aK꫎�h�����
�����e��]��}f���
2�e���	3oeD����H�o�d#�=Q�����+ɱN��jB4�E���t���b�]�2`������F���
�96}��Y"����V�H	�-|Ӊ�j�����v�
���"�kn9��X�d��.�/����|�i��H�S~��Y���l��>���ކ'#�*~K�&Z�R��-t���<�-��d��5�S��on�T_5	����7J�M�u��J�M\~p}:��e;o��!�	�p]n�f4���o�q�ꖯ�ѠJ�{P�ԣ��F0�dh=��2'Z<�>�X�`��C�uv�)�3L�&a,xx"g^S�bX{O)w~7�D-��#S8�s�H��6�:eMT&88����se�H?:q�*kov�Y
���me\�yG��+?�����B؟s�#�x��>�U���N�.�e��_s�ADYU�r'@O�}NT,���e%��e����%R5Z�w�f��^�Dr�T�n�]�
B��hȢ��������o��GL��������yl��%v��˾���w�*_����@�E��������K��j�;�A���%�6K��@�L���0V]I�&�1��s�ki��/c�i{&<���M��#u$1j0EE�X��y����<fX�4����>�׻��r����������72,M�S p����`w�wc�lfAy��&�����;n�U9�dn��L/*�T��;+h�l�Q@;��#�dQׅCJ�Ů����X�v\�EC�6��S9٫��I�p�d��yva���¶�L�@+*/��O!�1������+�P]]�ɉjG #�<�O��d�+���c� �E�GQ��hD���X���
�vZ��ad{��u�p>c�R[˗�Bw�8�[�MD6p���0�6_�=Pp]���J#@�����B3"b�	& ��ބڣ %O��k� j2���W�ԗh8�B� [����[.��_<���+����E �sݨ-��%���\��.��j=%�ű�_W� ��b�QU7V^uv�G�a�L��Z��A�ft���]����QقM3ς&ͺOS�5GǸ������������P=ge>�z�+.`O\Y6x���Y��/��w�6�eHH6���h5C�IP��@2'<o��t����c�f��s��>ւ�Y�o�ġ��Y��I|,4:��OS4����3h�oI�02���͢����)���i�sv!uԂ�{��UA2��x�L���>��ş5���e��7nSd���(a���ѻ<
�f�ۆf��V�X�-�Q�UTd��Z&E˱@��� \m�r�\=pׅC#���	�=�vH��q���Ґ=�?��+*�ux���)�2/��|�ޏ>�ܖ�L��X5L��>�3M����w�y�ne�}��a�Q����2�n`��Lu*�JT}��}�GRq7�ߣ��|z���*ò��p�jS@�D@�p��>$|S*�$$�޺�o�0c����t(ԅ��N�c����#�կ���XD�����
��,E�L	޽^��B��Q�g��Ҿp�����t#覲�bU�d}��[\C�z����a^�ܷ�Dn%�;�Y����G���7�	"���h ��w٠\׿�=9Ma�+�i?w�Y����X���ǳ9@�Az�-۫�m��+yx;����A
�QL���8wS�2�`!�uXU�lEb�������S �ȕ�"��ּ���>�0����x�ʛ)���<���Xe�B�O� ˗���X[�ݣ�E�Ɂ�5Ԅ�.�qV����/a���AV��ڏ� ��bQ;��=�{t���3]�U�.d��\:3OO��Y����,�t`IP�&5��Y�Qr�t^��`�������S�¾ S�-���JwYX=���1�MV^��(���F����K$r�˵W��pڠA�U$d��B]ISK���4�j19w�%���j��,й)��?�d��wu�V;퉴t��#&�i���YW�ŭ����A�{�o���5�FRl6��C��h�^p�\~�-��Z�N@���g�7�=�A3o��R*k�ԝ�x��`��,�\9��u؅���O��.���:S%�l7��?�i�7M�5��,����Mg"�%��xi ̅�5[�_���hiW�ԞIW���w������+Y���12j3	,ǳP�b�����Ma˲��'v�����Q�l���U�@�����;�M�c��g�b���[?P�{�x�0�R�ط7[���A"`��&>H��a�Y}��H�,0���s�	��^�^�=��O�򊵷R+YV�1� [BJκx��#e��JQrR���~m>���Os���Nr�3��)nF��6����ɊR���	�Ӽ��&