XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��� ����{YN�T�m��3�N>�Ch]�#*V�~��p44��TaJ["�9D�P=9GZ������ʹ1k�R {(g���M�_Ϋ����P=`3$^�)Q��]y��o���A�E�T�L�˶B�������~J��o�1�f��c�~�Fҟ���RG9�.����9�e�U��/�����GUy"�k�yV�	,�����>�QK�?O9�u.]j���;���_@�Qr:$�����Ɏ��F�i�; ���=����VɓE���|5{�¦�6�{'�KZ�zS�Lu6�4N'n�P�uW�����0�����$�_��F��Y��mu�-�."�
\�X��^�94�\.��,-t��?EdvBMM�V6W{H%�6�������(���/���j 9D�FU�T /�j�E�(��K]�����dXG�����f��H���@:E�⬢�+&;��OLBN�s�EYs���B}����/������ !�*���9E~)��/=2�4�k������+[��a�'�������d�n��5sA����
W�*���>��`E�)�Z�O����I�I����V����q�(R������%1��;wx�CdlƬ��f�IN�^�A`L���(� 3���uF_q����9 ��X6H�ʆ���m�&�ʦ�\��p��構��ů�י�m,��ܶ��}q�mw*3{���̞Ѭ�}�(2�d���[;�j>�·�Cω�"�Cj4��R\LF YBC7�XlxVHYEB    1421     7a0&�u,�&E���`�e���7�y�H��]y/��-�]�F;�-�(d�T=�)2�}��AeP
R�L�1[����=@{,c/] ���LYL���hB�cʙ����R�g�뽖$}ԛ�|�$8�V��Ⓐ(4F�@�aG1Q����i�p.��h�X"gl� �����*دw�z�Rs5��`0E���"�/��$��ӵ2���U*��>��,��۾��7�n�]>BLD�,fY�"<�O#�~°rvw'�f�Ś�,#�����q�?Bl���cj�E�(��6���e�+�OB]��Fg�q]�} ���9��f�vË����?O�E�d�a."j4��ª��lb��l,9]:�a;`�ܷ{&���m�3l��e�ܳ@Zyۼ�<JC((m���`O��-�/��kqh����7t}����<Z�ۺmBm���{����]��8����)o�,������b�i���=�n�pB�;�|PM����kS��b'���btDj�ø�=����F*שbT=��o_����)y݅�a�[I�ܛ�d/���f遢�_��+W�G�-���)�����iea&}ND�A��������.�ǚ5��dO|Gυ���y0�|��@MS=�f��Y�V�1{Sx�;�Zf��ۧ߾f��q���NT
Q�6��3�}R��|�&��C��/	��iYU����Ј|���W������Q�gI�|��)"ЇVHTP���;j6GqF�(K�0�S�F�W�w˘�X`'c��Wz��{��<�%B�����Nt�_҂ϹD��)^�wK�����c΀Vu,��z
�������������A�Z���5��GM(�t<0�{�B'�&\��SL�}f�F艴�
1B�&��F썾c��!�O� ��[P,�J���mǿO���qV?��qV�0�����N�yAP�a&��JV��9g#��n�;�8�"%o�)���*Q.�����Xq��H �o'���q��mp��� �}���uLU�ׇC�����KMC���\E��5�[�4+�}��N��Vk������EHǓ�g�L-��!Z�Ӟ
����p�K4�������xƆ:�gm�n�u� p��%%�zI��:F��-�[�C$�K�28�?�7(`I�*��o+�Y��»g܄.iɡ���׋-~����q�]�δ�E
��O�/ā�����#�� c�Pw�f�k�dB����"Vh^�Vٽx��Y�%)ZB�F �蕼�}&�F��I�	=�R�1��m�P&	aG��� 
�*�	<���p�N��1)KL��՜]�����:|�ϒ>r&؟�FG�:Y��yP��̜�	��r����7=w@��S�Ӝ�����[�[Pd���0!E�iKH�T��y��~�r�HLq'0#�B��wұ������8,��aԳ������� hl�ͦ��M7�+p ���(�
2b��5�u�8C�Ƣ�|h��]1�\�O�����黰�O䕶(?G�.JcKۙ �$'��e������bN!�?����^�_�n��22���#��|4�j�f{X�!P��$Q<X�KΕ-�V�j;����[���`=��y���J�<��s�y� _c�O^�GV��Ę�#9�{"��� �"�ɂ�E}��|ܟ#���~0]@����s�_.���4�#4�`���ւSM��\�Q1�:��y�'A���ѓ�����T�P� [�_����*=vS~��x�H���� ���{���tG�>�m���p݂���F�텏uߥ�qg�pk��� ���tﴺ��@��3����N$���]J�.+�|1� 4#��i&9�g��F@��S�eI��L�-�ڐR*���J~�zǨNPb��7�pdE������Ώ��-�8b�(�<=.������t��W