XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����ƛ�~L*��\m��"�*�6~
���q��{�R�^U2~��_�v���X�ݬּ��&I�j@ �[��u����T��YdB�����
����5L��:�22�l�mPtk~��T���^��D���XF"���K�������
"��>��J;�lXZ��qrY�ݬ���)��� ��r�T2����S{��
_�C���5Qf�asvO^��ͬw���N�YcH<fB�oD� ���{���79Q��^L7�6/�uH���(�P�	ŞEws�މZ��X�F2�涁8c�~p��ӯ�V>cD�"�k�ٟ�&�O�x!ltd�ӈ,mw� ��=�A�s�.��k��e7�>���1��Jd�QCT����V~��哅��m��L<��j��خ��[&�(��s�^��N��,����eP2>��d$� ��c�9`Z	N�꒝���q�?-[���c.�/]�Z�Lb�ʦ���KM�Q� �T*-z YCI[E��s�D�[vw��&j>c�ye,ُd^[�trt�ǘ��Ώ��8R���]�!�v����c��1f�ή��^\\�Y�4�k��nO��06��)����	a�kƍtD�!�3"O.G��p�{��u��tLt�(Kġ��f$J"^*r�:	A������qW�"Tr����E_��$�,���h��XI�]0�_YK�D����I�=�B9� ��Ѱ�S0a���b�Q�	��ͫ@�@�Q��ɕ��K�Y��L9���
;%O�2F\z6f�u�ϒ�s(��tXlxVHYEB    15bf     890�_4�������}�܇�f�,}�e�<���X˸�v��!T%\,CY��-��Sc{���{����K �������:�k{uzD���35\~s�	�wq���dM0bg��~(��I�A�h�ko�Ή����a(��J�/Y����I.GC�
˺g*?N�~
n���
'�尢
���Qqu�+���zf-�ϰ*�*n�j:A�$*�y�!��=�%/��j<�%�L2Ϛ��"P2L�Yv�{3d���ƹ.f(������q�]�8��	ٿ`U�kY<ND�14OӂG�0�㱹'DS&�ȑ6>�ժ������"2\�����th��u;�]�Z�'�([p�ip���+�_�l�����w�7l՞6'.�Jx��`oH�'U؟q(&���=R�ϥ�5">�|ԍD�^�h4����17�
��zb�[P��T�Y��WOr��% �S�@Ŝ��&V�4����	35��DBk�6z�f��=����1�N�̎�d�y��܀n����`��iݻ{.�Q36"PDzC/��iauZz@Ǌ�%:�1�q���VX���Z� �H���:��`ή�Pn�ͥ�ђ׿���6�r�O���P��$ۇLT���g@y��CϬ���Rj{�84�a65KL8�q�O-I�@�Oi1}|)/m Gb�*(��T������.�!qd.�)G�qx)~��Q�T�X�?�35�1�9O���Ea�}@
���X�f��P��o�q��Lo���&��Ke��J�}�)�`� bz�|���hK_wm�h�%�S��
�T@l���'M��?h8/����HzA�к��F?����V�!�=5�������
���N�7e	��QW���c����7�~�&Ӻ�$�X�s�n�}@7��6�[��b�d �o
_*31�ta�x8"����`M\&�Ҥ.��T���ɧ3�!���(���;����X][��	��S�+�lw�f4�=k��P��|����Fl�L��2[�����%��k	ّ�٨O4UK�LJ��޶�9��H<�V�����C�F�#]�r�˪�R�a������q�#� ���0��Ǌ����� ��J׾��N-ؓ�G�����\�t�\9P_������J��2mo`T�mv5WӚY��Q[���3�&�9�����(���R:���P�b��7o#�E��vw��=����4HT�m��|-+�<'���.�E�-�������^h�?��[4�3�у�d�'!��EQJ��#�Xᮯ3��s�5�v�.2��Vj�E���;H�c��.ٙ�<:K������$�Q��v��1��TU~���>��v���!�^����vVJ��E�1�0%�u6�B�n$�G����`��Ї$�j���tT��j"�tdq�^�(^4�i�W���TE�ۜB����g��8K�a�J��W;I�Gh��z 7��ƾ0Q����j��bd�?dr��ǣ
%��Kh���
���_jf�lB�ڀQWo�Z��;|H{`�o����a���2Lİm9�ҏ��a؏uܾ �z�Q?�����{��:�3����'�J*b�\v��>S�ϟ�KDt�AS=��ќ�x����q��X�ڂ�qt��A�P�������g�TR�PPQ�fӅp�e��x�pH��1���b�mLSau~�6ٶ}���<���8�UJi�Z��n�X%|fi�0��,4°D�N~��Z3��j8lKI��}��Wp� ��EHx)���2����	(�Q%7WP��fo՝��Kt�1u*��ϣ6lI���!��������Kd.hDk=�pY×��c���z�+m�iB�>��v���T�R�9�k�}�=�"������#����9���h�@]]�gZ$��y�.3.�D�����Tni;y���aɱdi���:6dLL�umpC�$җ��ʤe��9U�w��8��O�ǝ�*΋�s�&�w��8�UT�C�m[*��U��(a�`K,�K��Y��z�\��s�2���*u��k�*
� P���)��R��ADgeۭ�(�-&m�%, �GS��[\Cb�5�tGA��:�f'�,ًx5��v��� �6�h�����z�v��Ѝ��̴�1Å�K�H�k�d*�Ɨ�/|���F(�!sm�z