XlxV64EB    fa00    26d0�B�&�7WuPG���+�(��6�:9�8<C�!9%��r��3|Fu$AB���r	��e=o����U��ǵ���";1ˎ��F���֍Y��2�,��y+6mv�S�$i��dh����%Y�@���+q�U�N�} ��t�B|w���ֺ�	�G|Lu!�X�� #U��M���#[��Z X�u7q�	�ߘ��
�:!��w;��{}�٨?i�.�d.�l+�H�V3coX��z��v~�?�Rit��9��6�8����`9��6c�����������z��`�N��n5���n����ʋ���s&0ѵe�g�~!�~YՃ]�֞1&XZ5e0�������ߦ�Nc�%��&PV4�OEչ� kc4�f%܂�b�
���#�"��ÿ��A�_`K���$^W��ۢ���%`�lvax�wh�| ^N~��r|�<�P��.u�7�U�\�Wdg2G�fc�g6�4ey벒���]��~� �+�x@g���hh;U��RƆ�|]S�Y���\1�##����QRW�&�Z��C�����~W�υ��sl�W���_��\YET������yhB�o���P���Fy۲C�9�a��2��������{�t���7�RpY�������!O8�We6_�����q�1�e�R�IJmK��wv͎�q/���b�8� R���v�_��`}��S��*.a�f}�uxP�!�Y�=TT�U��!u}�=VS���=5/�*ͷ�k��[����w�;a0�xq���r�������"�������Ϸ�2���\��XP3�Jcuߗ��Ϣ)��(�#8"��+e�dZݬT�1a��Bt�|Y�҅��TuvίG�C�\":Jپ�9Gp9F8z��iȼ7�-�0���}C��ւ?����"�)��P$�-;D@D�����peC����l�^�ܘIJ�c�C�-NI�:+7i��?�� ��ދ��t�~ͅ&����z�oX�/,�����Ri�{Z���� �r��v
�m��ԕw��>j����s��)X���D]��)�7�a�H�3��O}�Aљ�pM}�3�����0|o��[��9��C����bO�E>���5̐�Ң�B�tR�0�Q�N]'ѱ������k�
�&�����b����ua$4��y)	H�5[Q)+���}�j�<I���ʱK*�u��A\4�~�j
9��S�v�����+%[-	�W'��pXd�ĉg����C��p�NTjXPa���G-�&�#Y�J��GҞ&��^��I�3� =�j�_�-C��	h����I�U�[q����q]�5E5q����0/\��D����k����Q��0^^��gM�]���o�p!Γ��r<��0cCZ���~���P5����sA2���=.����T'P'���A��.�(��l~��L�E?1n4�ܜ�����-�C���/�,�Є��b�,Ͳ4�gP>6ηM6�Q����Y�(p��뉔�|BDo/�Ӵ����#ս'�v�x�;֫ef�N�?�K�Т-��-�Wb�k,{���٨���O�3(|
RH0�M_��8���V�����"^�: ����#rݍՀ'q�(\���{"$��SE_:r��T#[���SZ�v9�t�,6�؋.iT��K��ܟuSY�	��5�D����|��t�$0d��eh��o�:h��%�5W 6�%�WP?����6�P���7�I�z�P�)�.�2-Rby/֌�]��/�wع�S<���=N�ώ'�h�t" �!<�c�%�_�MI���p0+6Y����I�:�5%48:rV-�/����h�4A�(.(� c�!>4/��J�3&K��K
]�r-S��R:�^(�匥��#�V'��\�0�Oʦ��x�7�( {��[��}I�Ƨ�V�=���3�ػI\���;Š�V��:@0҆�X�����ZM�R���HZ�9��<��ߙl�k�f�a ;�
����j��tL����{�bP����H�3k��,%dPڎ�},�ٻZ��ǈ9#c|M�ԏO��$�)Biwtߩ����,��H���~x��c^a�������8��ub9ܟx_p�����dw���G,�ʓ���8In���������ͷ���NC{M�r��?7b�P�~aX�i9~��㲅�o�����k��a����x`�DE�-�>u��'��<�.H��F\�iy�!V'H#kdV��
���u��o�b�ۥO$�lA�8�c�R�'Y�j�x�cT4��S�/�����#��D�����R��gQMӑ.7���4�]M����$�E}
~��5��=�8r�?��XN�C~i��T�)�����������QD٧k���c�{�m�ˍ�p�L�o��!�H�9]j��f��[�ga�����fh��EIg���9��8\q������!�*j�\-��r�8�`g"��h�(�d_����v�����.�X�X��*. O�u~H�78�zD�������9�q ]2+7Jb�ޫj���6,K}�@�3#񬮯�Ɋ(o�`���Y�T��K�][�띶v��N�Ȕ>�	������3%\�cB�0U�@�>�Ag�c��:��`q	��$7"�J��j���4���W��j��OZ+�PNa�կ�:r��KE��e⤆|{A���� ]e�`����x��;!���W�,d�?���Aw����,�q*K�� YM^Š;�ޗ�l^k�[ŽO��}{�+x^��SSBS1�D�E�o�H4�<hFKwJ#Դ��B3�z���
ߋ�	��}%�*zWE�TY��:���q�d�W�
]zEsz��^,"æn	����r�G',�f�?`� E
��,�4i@�����఻/�w�b�C�A0���W���
a�S���T��X�X��?(yG��f�1�w:���DMóeS1f�����g`!0�{����}��x�)�)²��"ņv��;���t������Q��;�n��^R�WG����iI
����G���ρ�:������	&f�J��iL�jHI��Gn1cNSܫ�$V�l�&�Z��T�H>�DK�
j.�(A���I�b%%M���u���p�����FH<5����i�B��~D�q�9g=�1��V��/!���oZ����ޓ`1���DF� }�G��q�Å�7�.pd"���rk�.������/�Ig��K|<~�Z��l��0(�psX�=�ZʾY�ſ�v�/]{�4�@Z�ZJ�H�x-�þ��(u
�A�2ת2L<��B��b3� �zت�����eQ����7j"����A�P2�㪡a<]o�
�
�fZC��mg��<�
��n~��q
Mn۞A��8���$cpW���H��u�p��l�����Y-���z������e �f�
�;#:���8�3}8���%+ǻ㛶A��. ƅ7��,]����X�b�gC��C��<�fj�a������زo-�{�#���b8�r�Ñ�@U�R����B�P�c�w�|�\A�Z���B�q`2��%W��[Mp4��-�����%�b�r��4>���^>�Zؒh�S!�����d`U� {i��A�<�`�mhP��p���O�ئ�g���a4V����qY�>���Y�ܻ106�	S}(��9Gs�ᶃL|:�^_�*7�l�M�i��\�h؜�T}��\Pz�ez�$ي�\�[
:;Že���0ĉ*��5R8����&��B݋��8��f��$Qe�u��K�^�?D*\b�{B��25�)a���7�`�e�nj@�86h90�,d�2{ JG��"��|��V��&��9`������$]|S;1a�� D�Ϛ�ت�-4�֚Y��-%ߠ��ȏ�|9o���[�بf	Q=ӻ���>;�2�_7L�X�Σ���SLk3Xt�3� �����tz��f���7�9몜0�6����� ��0x�\�81�H9������h�/���a��ڑ
V'��m/����=N��E��A��D�)��~6�_}V�%���*+
 "ӧ����Էv��<ƴ�u�o8>��$��\~�`TrҝP�,�I����O+o�am�)NG�	&(�X�)帠*���3D�©-܀��!��̙
��sl%�2�:~k�v`�Y�f,Vȟ�EU^ya��a�L��T�]*a�xzG��_��iD��Ch���g���8��\?�^�x���(�v0��>�A#���R��![P�b�ە %��r�M2}�tW�Ռ���֟ u�8Ȩv+�������-ˏH��6��K��e��m7���CaR��?Pn�Q=Q�u9&��a�au�}��d*m��? Zi�^h3����5o��M1��Z?y���7d�p��Ԗ�Ɔ��9�	W�ufX��-gNnN�2G��ṗjk�GZ�P��k�t���0��а�?ޕ;�d��V����}���E?�M5�A�k��l�	Pj/y�B\1��?�"Hy�{W�q.��ˊ�f,��*���i<,�Ń��1?�V�%���J>�B�^��'��x�(��;�������छ����.Re�����*���u?k�;Di�LR�P��S|>y�{�|y�����2�@u��äo�b�����w��M�̬/R���Ņ|���L�Al��o��}%�\�;��6xMq���ù�`>�P�����x��Ͳ�@Q�5u�����I�Gd�t�'�g΁o���b�W�6�4!Hܝ�3ڻ���Z�����W�h:��ш�n�Vr�?��[�
���X��Y�5�"�3-��Cv���̣�nVW�7����
_�r���d���i&�"5n5�Hڅ~!Y�āM:�ۦ)3�d��� �.��k�����]�̫�$����0�X7�;���^�\�E���L�i5���=?�I\|�I���$���Xidѭ�q�
z�KJq�'�+��,�y�,ܘx���J\���p<�}��Q�
?.W��O��p	�S������h��#U`X6(V[}`�=���z��銷��F�#s����B9����،�X��)>�-X�m@*��V]>���_Q����Z6�u\<f֠�g@�
s��6��G���9ʓ��='��^$u�a7:�K�Ar�q����CTf6�X��Ʒx] FHzt��)�п`vX��Iޏ���4�A�$͈��q͑�.E��R�^Y���z�${;�}�	�L�� ��U��M�ǈ[:D�W�ۑ��$a)��W1�<�y?.�������,��r9h�~u~^z�9����t��_���~6�L��u�``M�� 0F�V�8�	i0#bтin7��,�����	�~h�%�����
�0ƶ�3@E_<`�*{\��W!�Z��'�.�qk�q�Ǚw{1K���|�r\�q��ʥ"pNY���;_�̆�\�0]�Q�}�X�Q�;�:���W�e\��7�Ƶ����-N�|%��)L�`N��.V�s;E�&@\�F��"�kb[�� p~�X�#�.q��W�'u�j_$�r [j���O��qj�g�L�{�m���F2:�.��o±|
�!��^�\�;��ub���
{%��۶�
���j���F�l��"k5+���C���!E ^�R��K�[9�"�e��%���]D�VJ�C���E%���|���@x�N~���z�EOA̗>���L�Mğ���S���s+�t��x�N �K/�8��U�ְ��t���j;ұ	��@��'	�^q��kgP_��gŠ�K{5�-r�D�4��ȡ�V#�UۇU
Zxɥ��T�wN��b��bfCI8���Z�ݦ\���Y<{��KF�&f߿�C�`�ê����H��Pn����#V��
��/�_�^�v1�ƻ#=�^�M�LQ����|Vt�W�#���Â-o���SgW�a��d�]��y�5�@L �64�vj��Ǹo�3�*�K�W����Y�y}�G�8��U����U~�*�a�|��TIr�S�m9���Bd������ڢ�u���m�"e'�L�����L�zП �褁_��vk_ʭ�����|� ӫ�J�2?d���"��,~;s�1�2���PShٞWO=���lɵ���@.�ҟ������]��T}���C����&�[^a\�������T���DISc�G`�ph��&�]on���"���]ل��ө�xZ�����l��,�w����T�٩pm1m�/�����/-q�_��i�{<5�_n,�i�L�n�u����%�YMk����˵i�H�����ÌP��p�w�0)AOsX�a�4��'%@wTQ
��~M���EA�� ��K��dHzx5�\�H"U���\���B	�_&g�M�6�{C4��x��y�l�%O1���q���Z�����I�9�
�P �݃{&K����za����)�������x��Y�*�Y}R�l+aP=���b�s%	���S���|�K�ò�O����-�����*�mڅ��ѿ����p��ꙁ"�@p&w�;Ցx�+
FW��%���/�U��y�$`V�M@_U檢������tjҕB,I�T�7J,l�twI�F�$$ډ��鳹�:ԹEF!�Y�L��oYN�R���Kl��P <T^w�����������ɧ�UtD��^���I2��S:w��ǯ@�9�`t��[�2�>TY"�C����9M*�R�b��6���]K�����ç���}"�r�K�]y&��.� ^���rkr���bUa$Fg�@T��*���s��q�&�̬gE~��Dl�ASd�l���p�TC���.j�˂`hs݆ů8$&��#;�,�N-�7ۼ�db󮱕�p#}~j�,BU�[>��8�k��U�����q$�bR.�H�@ĞYU@�;lN��B���;3	��]�z��H{)8��TU�1���ҵÅ9��O^&��=��6�3�G��&4��E]�uS�>�X2��#��[x:�-w4+��Oи؎��e��ˬ v�Mj����	��Z�֒�ȫ�V��ٟ%0�1�N^z�\y��؏��)�
yA�>v���0�T�'�|�re�V�H�SӀ�� ���Dq�\��p}
�t@b9�#��ئ>W��X�K�L��ə���%]A�l"${��\͓�0�hnU<	��F��:Im���
[�C�J��X�0f��P����!4�O��v���w"�3��B��-����o��4ߺ�/kҳ��u�vz�����ؓ�g�8����7�:V�<Aa83>e�KW֪��k�c��	?	�)䒹8�=&t�P�m�Tw�,5�1���&�HQ��J�y� ��ٱ�����5)ޱY+by�!�
DnkNwN�y�~9���לj��34��:1hуP�?�bN#�c9ou���X���{�A�Pz��A[a�\���J��
`�k��V�O͸]�y��s�~�Z ��z�F��a�[�=��œM,������e.0@�R�{z�I}7�U�-J�7���EF��Ĳ�?����$��3�Ok��p�/��ݙ���8>o���RY�5�����\�5.�G��@^�����D�.�������ԩs:�D.��9�۽�e����̸(�\�A_)(~�9ăD/����Hq�����7DP
��?Y��ɫ:i���UT�:�kP���${"�6�ٚ����Ax���/�g��2'/U��?���v�;���?^c�1�,%�e��y��U��?�$�)�n<c�4��6��.b��Yh<�>���1�~����/+��b�")g��d
�8����˃��`�; a�{�/d� ��h8ʳ6)�@����%5 �ˬ�^y�g����l�	L�ntB����Q &��U��GEa�LNB#��**W��W a���A�|dXB�#&�}b�h���7iݨ
�qd0a�gy�pvPN7?�����%�K*R�:�'�W2�ӳ�`LV������u�p���B72� ɻgu��̉d\n��������ګBo�٩�{�t=�u� ���rJ�h�q�W'�SH[ݘ��pTAJ͈�l��>�bO����d��,u#S��ox��jԮ�,�������w4��2�-��T*�/�f���ΘD�?���������!B?�UQ%��$ㆹ]S��eZ;�U�4sT$��3o��*b��8v�|-,h�Y�葱�pp�x93��?r[�����ƶ��l���B:�nq��ؘ�]7��������4~y������$WJ@�U��h��#�!x�"�9 1�3Z��
PP����j��cb��`΄�J�cC��g�gV�]�c�:>�-{���@A��n����`�[E�&�w�FS�'/��l��.̾͛Tj��j[�`��������;/_�VQ5�3z/���#��c��#t�y �����O��&EU�>������4#!���[�g1n�]LCd6�g[��+��I��੄Y�Eu�*�9���!ޠ�'����I��wA�����M�v���)<Uud�xw��{��X��P�XIlsU���-s�DJe��7B�͠�oQ����@�A�z���\e��  ����e����c ��ظ���j�͈���h�%c2)j�	�y��}�NL˅�	��{z�;�?'-88ue��@4�=�Ssn�:�o�'����Z��r�|>��c�y9U����a�hKv�/�f�n�0"�dcQ��̷�XZ�~��ԋ�VJV��J�,S� ���D�~����-��� �ql��M�&%�!SD;Ro�V�X_�~�-�9Ď�9�\ؗG��f���*�vY���cfr��Q�-׋~8d�>�L�B3H�"_:wJ���~�����hl�FמG�/^��#c�z�]ӧ���߰������Dz��֏3k�|`8t������V�*�1st�G��(h��7A�8����Tx"�ly��.��!2Ml~ƲR��^�J��{�D_��2�|�������9���h0����VZ�Z����R6��A̛JP1����T��K�R�Ә�>f��0\�ۚ�?��{�0���'��dj7[�fR�b�V\p�_���[�ٜK�5p���x�G+�Ԛ�C긣�Px6��$��=�k�׉FD���,�����l<q{�cp�ل!��zv��\);����]T
a�����4�a�8_&=b�7`�u�D��^�b�E�g�v$62�h$]A��I@�_�8���O�,�zd���vK!�$��gY�� &:�d�Y��'��^���N4�H�D�%���f�B�F7��(�l�ô-�T��	.���X�EJc�#�R|��5� 3 ڧ�K��+��\�AM#�kY�2���0(�&_��_C���~~�������d*�7U��Wr� �CcS�v�������=�3�=99�k1�w�@k���*�����l/��j��	�v}	o;iR��u�n��P��*P'������?I�����li��x�wa����9N����QF\�Q�Ի/
����v���p��Ѣ�6$8�G�ӵ�;�r��V7N�8��ϫ�lS-�s�v1nF+R��ZKk�s�/Wي��q�Ӈ�&��oSq��y~{�1�dd��� �E(0�F0o.�I����+i��O��R�AbL�Ȋ��b��(7y�{�7)�%f����w�:��!<�gz=��]77�JR�]�_$-P^�����㌣��ze�z	/|IP�@鱧q5�B~`��|#�� ���ŭ�y��,���M^AM��~7�g(�^��_�V�XlxV64EB    7c6e    1440^�t��)cpAd�Q*� )�g$}u�!͒���|��<���5Q%W�W�9��C�w���I�����/�^�����jŠK�w����lYk��K�ۇf�5tW0A�;M�������a��H�vD���t���=���/8�nT���� �:7�z�~����\XN �t�j;H��׊�c��1R#���W����7�i-����D������1`��|��@xtB��7	��q�G 7M���m��"��5/U[�@�m���q6m�lr$�E�n:
�����Ej>	,o(��r�#����\�L*KV_��=皣%-^��Ⲿ�@]��`��"96a��\4�(8�C�Q1Q)��{��T�( �*�9챶EL	�{̖,���T�FhH9�^l�#U���ȵ�|����>֫�T��o⾡aڧX��Xc3���_'�gI�ͤQ�[k�Pdi�(k�3�cDoQq;I"7q����1�lr[E�G!�:H�#�Q�O�bÒQsO� �F��C곙R��J2fA��<=�`B4�`��B8�����-�飐>��c�����x���.Nһ�[ޒ�-�ј˖��ر�ivt.脭�aT N��E����	�"���pau�n�>��E���:����?�����oHYX���q+���msof��:@u�+ܠ
�Lϵ�(�"@
UcK�yX�W�ZL���gF_k
IV��#�Q{A KC��rZ�.���7����o�
JqG�<-M�K:na!x��n���P"l�&� fL.��4'#�j��
�º/��ʧ�l�풻K/��i��˙$[-�w|	:��
�N�@���^!����GY���-�(��ҀtC�t9�ho\@��%��K�n�wTDǈ�<жN޶"��^: ��ܝ������=}qe3c�|���'����
��]g�ӓp���`~�ܣ[�D(�%���*A9�e��!`Q��y���F(S�W��.0��j)�&�,]*��η�f{)��f��]���h�w�lΆ�V������4j���,���[�5�`E���G���W䰨'�;�	����"T��K&,��.7h/#1��>ᛟ�n�Z�)Z� �Ʒ�ƠM��qqA:N0?������������H�Yt�G�h��/�&�DZ�1Ј���Z""v�=z�!%��V��>aU=��a<o��.qғ��J����X+�&��	�|�zڞ�\�m�V��Y���x�#�8Pӂ����)���WBI�r#��^��Uh§��Q�5�
���[�3W��X{�;�nܙ>'��9h+|ޓø�|	�B�6A|T�Bn�z%��A�xM�di��S��;���F�g�UerB&�����a�:��+��<�Yy۲��
�2�&=O$�>�"s�0�{bJ��m6
t��GRBt&8s�B<��ȁ���������_�$��y�0�Z���z��9�؃�&?�4��<Oү-D"�����ܺ�G�\?NHa�	��&]pd���O�EHM� �\
o�ҎqBW"���h>�ߘ��_���N�ŵ�#�	N�[ô��'�P���9ql�o�`>o���#S�!=�,��Mv����'آܸ�RT��v䬇_�J���[����� �9��v�� �E��pt9��%/�,��kQ��	n�am��a��k�l5O�|���`�-C_��i��ڧbd�$P��`7c
e7^˔a/�LƬCK;�+�G�뙰���&�5���_�:S!�9��s��2L<1�鿲I����\r�N�g�9M��[Z~�f�������.<��%N��l��eu��� ������+Q�S��V��ފ90I^�_!�ᩦ����C�5$OS�-�u�b�l��n�=��t���9�,�_"���~�-��4AÎE�d�_�����}��$�	��i-E�b��7�o�S;w�bj�׻4�5R�^�{���d8���e5��
I�Nｯ�c�����LF�x�Y�ۘ��b-)Y m.y�S=�:8 ZM�]?.�Ŝk_}A*4m�^$��T{�����/9�a�@��'{:J�b�(�P�u�E6���-��I��{r��Bm8���Z�./�n�]H�xC�:�����|T��ķt�e��hr
��!�pb^�c��c
b0�HZ2�e�/�޹��85ƽ�t��^�~��ڍ�~3��?d�E�Б_����z�آ>��)�}9#)���qĦD�oy�&H�:4بrCƫ�i,���.=��#O���n6'@e��/6"�Y�b:�k�����p���k�����q��-��"T�i�攱\��d��Q�T��u�5۝��NvmFԿy9�OGܚ2DȬ�4���j�R�P9�`��A@��7�S������B��5g&+U�T��H:�ks����lb�}zՀ�j�`6b2��ͫV� �,��&>��$�0=ۉL��v'B Ds���*�JNZ��_���b����0B�l2-�\���uBO6G�*kI��6�8�ٓ�1iz���	#�����<�ɋ������ҋ�h(���}��{��(���lN+��%����Ss��I���I4U���D�96��$E�)�׎"�kNkD�9���9�̽�=��}�C8j���Q����)��,y�u]��%!s@7�>�<%�A��I�l��G�V����H�����T���#D�gI��:����#�)�yr�#3���-�̶Tj4�m��}���`�%�!n�d��Ƕ��e\+A����&�苘�����L�b��pR���c�@�K��4��*���Z�{�ڲeI00��P�M�9�&v�<
���75��W.)J��+z�"�ϙ匓���њ�{;��p��,���D�ӡ6�Q݌~�j�� l�Ñ��y���ԭAp'0Y�J��P[ "�V�U���Q_��o�
vm��������*¿�
6xcЬU���ܯS�x��f�q��(�b��/��g�|����|V�@�cA �>N���l;_l��/��rj���APGy[P=Y����<4(��Z켱	�Wf��Xfׂ~�_݁Y�%���X}&�����M�xRd��G�ADđɗ�}��'�����tL9Um���H���b �I,@�d2]�zs�t켞��*��Զ��#�����Qh����<���0���G�0Jk��n�wqH�#�N���ed��<'z�"�Djf�Y��E�����Ҿc,
"w>���� �v���/a���a�
2v�۽����A9���]�-�<��&}V�"/`*�r9
�tbM�fM뀬�~���9���1�FU &�"�:�Fn��j1!���}ٷ�;YW\N���!x�Fkպ-�3��\��|f�T<�+ s�l1kd��l�c=�E��]����/�fɑA0���l2$ݭLnM=lK��nF/����l�����aܓ�>b;k��Od��'.E��a!C��Pd���Mki�p�����b���	�&VsV*�����&&{�T5F�A�g�4�QL����vh��؆���5��jgh8�A��I*�a�)�/G���B�, �Ľ��ߗ6�O�������dR��t��cqv��w�wV��N�TQ���š��U���%�ή;d^�.��6��&f��p|��7jKaj�2���ք`V2}�]due�k�k\��+r���Ϊ��e�W�_]vj`� @�����8Ǹ����tV;��"2~�B��x��(�b�/��B�������ǆ�۳��j��2G��҅I��K����5��wh �(�o��8��W_�76r������enz�9�A�#���D��\U�}o)dH`��R޷�Ȓ����[+0	@̅6a���|�F�綰Vg��t3|Kﺈ�6|'*��TT�Pa�vʨ���k���(�)�jDq�c�����l�<��43��K����s[��g��qDln��u��1�R��y0��0FI�Lɂ>F�#�m��>��'ض$�����<Y��;b�\n�����i�a��Hc%H�m��bT��~9��j�� }&��</!�g(��t����=��Y�v7�_;r4�.��p4�:�*�'ЌZ�}�JPʲ�&2K W2��잗�E�().}��5��v�d��E�h�Rz����ٚ*�;�N��xO��meq#dAyPZw|i`���-ݳ2mW\�p�>x��A��x�?2b�ԡ}���s�4��X�ܔk��s����h�4��+��c$���T㧓��s��z$�}U��$� �-��()����y�1��L�m��EJ���X}�C�}���(<�� ��X0�7Tw`����ǳ?��Rm��Չ�;L[Nݷ+B\ w�E� /n�������d�)�aWPB�C�h].2h�>�z��5�ɡѨ�����l�d&����EEV�yT��L��N�������D�ke9j�<"����TT���=���7i�\�:�3��O�o��i4�a�; �0B���r�M��n$�d
��m�h�d��\hV�?�9u)j����a�:r�QKa/A	�)�S`��E*��J��wAf�+.^]��c���֤�B�_�W�u��<���A���E>BĮO1#/J��f�o��R|};��$�6
v_����7�B����S�Os`8�*��;7�N6�X�M�J�"�Ɔ"�wu.�;�n^�ej���87��w�|q��N�_��=�fP5_�B���L�A45R\|���zx`���iG�TH���<'�Gٻ�cyE��j�r�ר����-�m�dڇ�����?�#X�ȇD�6�D��IoQpM"'NSזF�3�!�m��@�N�ǐ5*8"�^)�tH%��cXAE��Go_;k�Zaq�1�	[���]�롅j��;���сbr�翹-@�6YMb
C>�Rt�S���v./fSW?5��9��r@&8X�����&�.g!��1s�< Z)�e'zX���Pc�|8�T���ݳ �f����lc�X�SO�π���!�Y����"pU�����}����uucgK�����1]�Ƚb��F� �kѸ��kle#S��ĕ=��q�V���!e�SQ�,!EmZ�YO�8l�!��Ȟ�h�/
N����Ju���h͓��
̋>�_u�����