XlxV64EB     e06     690 m�50���=�_�r�F{F�/B
���hHb�r�i`���X'�'%���NZ�OP�L�-5�����&�����"��A����B��2�೽�gt�%L�F���9x���[<�~��U��DT�2 �%V��[��+��䕰�����4��໳$� �����Dt�+�&����ި'��hsH��R�I�m�B�'@��5�Ƙ���7���B^@�������=n3�����ӗ��;x��D��y8B|���y�:�}��x�7�k�&�!x!�'m�5��X�~��)$H���sM˥�p@#����-�n�]�nxC<��@��p����;��9Mt���l㡣Cu�4�{�i2Z��ڧ<I	)�$V��+o���!����X�K�G<$]�(1��|�z9���� �ޕ"^E�9�Q���_&oD\Bv��t�ɊTOq	��;Y�2m��[ɛ鉅�x�_�S�a�!EǮsc�ڭ��A츙�;W��r�Y���5����3^�V��`|Ձ���Y�K�,��3�'�3D��ط^��/�5'� GG���u��b1�w/+]���*��r���/��+�}󌭻'���դ�TɁ��������i����j��p��%�b���B^s=݄>q�.��������֝鮖��h/�R�:�b;���N�@�Q�o	�)�;_���3��)t���ˏ�Lʺ
" �?�[�uxi�y�.��ͷp��[�U(j���\��@���꒘$�޷a��I��X?vi�Ruc����bL�z��Ǝ5	gO �$�)�M�VOg� ����?|�S�;A�(Us�	��W�x�]��l��l��^����R���wϖ�����|����6���%��v��%�Ę2Q��^m��=�((O'�>�1����9��m+T�*���lX�"K���]��(�r�:�'�����#��eJ���oc.�'��K�S�[�fZƦ`��>u�!tX����#�S?�O�:�1�]ǅ6��O|��KW1���&�����J�thEq)L���xM�(�h���O��(���Y�w��hQ�4B!
��J�n��d2�����R��t��{�T���)i������譊_��i;<'�*���G>,z`?R<���㵆V�ބ�/&A:���`����%���F������$�(�5��@yo ��;L�\b#2��u6@Xh����*G[���::Ŋ�.�1�/|V];Q�)Z
�<�"6�+H��{-��1�
Ӕ�'�d�AK;�O�̍�&Q(�7#��
��`�gĉL~���V��RvA!����pQ���[�9�*m(�����[~��DjU{��Z
~��!��8�Ϡ+��x��xNa�7�P�Eg���_Z���HNu�ߌ�q+���3H3��Z>E�Dn0�8N0��[���l>p��8Srl+=]���/�z<Ӫ��e�g���J��$�`�ٻ��p�j�?�)����Ym6=��sse��I�ĘJ�����oò�s���yA��w�+Pɬ�+�)V�<�n4����ƛ�]#N	@1z?�-}���+a��s{o�<!0�Ҍ��HZM�cְ`!|�I"|kL�Z���_t��)��(���-�+�뙥ǀz����$s�3���,W'