XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��GtK�v���B�8�;P�ާ;�#떄ɀ	�7�:��/��vn��PT����8������J
ZZ%�z0y�7fH�D��0�u��qK�� �>����Ai�;���'aA{���>N�O)�W�1y�=�2�]��-��>��7zf��3��֬�1�B���	��!�EW7&iG_$Ԯ�w�%��n6J��1]^��=�O�bw���d�Y�O��K�r#���
��T��f�|ا_�bWoB�*��3.�Kȯ��E�"9�b�����k=��D�U��Ď)h��f*���&����D�
!}����M�Q.����<1�OSg���T/�4�8ӣ�yc�+Ȧ ���"0�+#^Tu�c�txX��<�]��4l@�qO��\G]�(ta�"P�e�JF1�F$´�[�������Bmc�e�����>V�S�`.�?L���h�rd'T�)	<�7�m�B�����^�����,����U�Q�p�he//C��Z��r��o4��d .%�d�'��w�:����>�&��c�:�+P1����fl�z����2O�����L �r��>�ld�̅���e����n�M6�~ �3+{e�u-��o��yu���(�J0|喦A����^��I�|�����x��u��4V� ��_�~�"T�cn����q&۬���`IYg:�d�2kk���X^��A����J;y;��k[̤%���O/Kwwe,n��=�g��y���u�g:G�XlxVHYEB    3da6     fb0��j�k�ݗ����{�a
vR����
����9!�%�,xi��^����>���U�y�P��f�8�:UO�wd�J�:X�
݅Q�� F�A�~�@�nѕB9�z�T���S;ft�@��¸�E8v�)���>�D_�?��݀⠱:�C��l��k���TT�m�|&�J����66'9���4����]s7?j�܅!2�K��Ż~���z}�A���P�q�ĸ�6Z��L���ͩ���Y�G���N[�e���fSob���k�`I��~-y�B�	dz��+���x��pӁH�R��"�T��b�a���K'�_�-�zf�m����:�, �T.�n �
�"RĿ.��R�9�����㐬�#�o��T���$�Z�zf�DSS淺m�������W/���v��,Y�{l��7XE\���Ɵ>��S_wo i 5�R��/���/�2��(�?c�10�p�!T����F�GR�����sl�M�(�����y����E�9FyU��,�M��ӧ�@��ƚk������CD���}�3]]��� ��k�Ō�cs���ꂫ�9;�������"]�́��`��^=ݱ������ئ�)�єm>��
ny@E��;����#�$Ss?;�7��Q�>o6�4�эh1��#��?��_�Jj�ca�XF�R�y��8�f��9}�uN���*�dVc�1Wk���{�s���ݨl�1$���~fߔ�
ڿ���_O+}]�x�@�&����L� (����v�`��lX�࿨�K�r��Z;��K-��8���7�U'o!��6�\���Ö���P�?L*������f��R���]�O���c}���H R+���:
t�]D&��d����y6G��}2-(���6M��B�\uM�����T�J��C^\�:"6ܶ^����)�U0�)V|�������t��|]g܂����'�����)�@�ց�(�Q���n{�YW�\z��(�{�����w%m���W�^���F���A�TF�[m'�՞�&q{�)+W������]C�~�d3�F�,g�1(��?��>��K�5�Y	9�q���]�=րcu@���W�v�� �)���+�5�������K��sڻ�S(1�L�9�t��(�u=ǆ�
����iRk���ǃ�z�&¬|�
��xzCg���E�#C6?;XۤS�nxB����E��Ztr�xu����bs �E����U���2� �0�����W!�<��{�V�p�YHX��M�Z��}��u�N�&v�{�l�w��m���r�Zo�p�=k�kW����R� 
�E�i��?�(�����s�ԶB�T����/��8�>.��򜕽,lY�B��݀Q�(]���C��1���d��5�L��l�jhcAi�K="�QM�����ώ/n��>g�W���P�8�'���z�N��V��n�#���P6�\�?����
@�+��wj�GX���\�x��:9��x�+���_�'�v������q�{�s	�YP��E��y�IB�X�)�ɩ㡤C����"�U;~��8w��������S�z�'j ���6:���o�ۍ'L�1���{i���D�C�9*eos������=�	�P�T]K�k�k�����ÖJY�"�P!#k���*��I���P���kҊ��G)
�Z7��Om�vf��c�l�����@A���ڂ!M�r��)<��Όs��W�����{Bb;�:v���xs�~����Xk�E�~�߅��f҇��T�Fv.�&��g�;8�ݟ�N�J=q����]�,���f��@����Ceμ���[5WD�x�תaK��x����@n���b�万BD\�?ajW�?�d-���$V��x�o�v���.bz�Q �LȗQ�^��9u�ݔ��ơ�Z+�v^�!�������yw�_zpޜ�S	��p(Z:���<�͎{�>R6�TE��1�y�P�8�aë�@��H�XZ�]ۉl���Vc ���j8�������k�P|-���W�(2��z��m��ļRo?�7P������=����?�b�Ńt�X�R�G�Tz!�1��h��B/R�3�n[OcԶ���Rbaݧ\�U�*>�3x�h�j��qD�!_��\<#������J���8_	�{9;�7Dk�W��.�Y�5�"C=�2����_"�s���GB���1㴬�y�׎+�	�2Z����@�
>^�̪Ӄ��4,�>7��2�<v���g[�[S@d���j�9gÒe���e!���;+C���3A�+b��u(����}����mR�pM����<�2�KX|T��fH& <ݎS���;!]��3E��6��y���L��EXU֜��~��q�8����X.�����d�{ �MgBx����.�(h��dZ�?w#�|�,�.��"+Oa�{�B�=O7h:�����	����s..��s8��( ��_�+1?�����4���[_��5��|B]ϧ�OբH�O���%3r��G���jw����2���D&�&5
���K��̶+�Q�I��ߠL^�+�|��v�1{<@xg��ʚ�iÏTpK����/t�����2�X�d����u)W;��׋\�b��P:$���\Ǚ��-}㾆[]Ǵ�ꈿ�.�1�e/<a��ND��/
��n�-[��׍Q:k���r� ;Ԯ�q�q�����&��|����-$���Cq*�g�I��ԛ�t������5<0�����| b~a��,J��Ni�wJ~��-&o���������ڦd����TT]����O�w%I���I0�B 0��������j> ���vxM-zL�MF�&�2�ہ-b�V�� Ѷ֢?�QA�w��~�T���w�S|'[~�\��Z��`<6���V_n
4`���m����b�`��V �!?�\�ZLC`�8˯���9���H��6�"����Z�����?B����(2���`�VM�C3���L�H���w�S��#�վ�ۯ���+�l*S��x���q7(R�y��w�� CT{�Q`�X�|��[��W�@�6�Z�=�>J���	u�?��3O��8V�ZO+�rk�as�1}�">�W�(ߪ wƼ
�E�����\/s�}�J��QQ,��B/�	=�aƹ������o�-n^hXvz ��M��ˇ���� ��盂Bri��ә��}���&�S��S�m�L�w��A���C�uMw�V7����5w֧yG�`�Գ��3��s6�N~�Q�[5��g�;�Ox9�A��������X�h�bE�v|�>��jG��	K�m��g@��%�m�*KX��xю�	�W+J�A���~|߼l�/�(�|a�bZ� ���6J렫�2�zm9��I�P��+��Ѓ��EWK��$H2'��S`�}�b�F�������%�jV��`�-cٹ����Ի���������U�|Y�Mp�8J��T�M�߳�ïTj�	�m�e]�����=Se~@6�ap\��VX���	
،sc���<�#]����p�Yx��->%�g��*<P{�ϥa u*��q\��MIҥq�K@��D�H��ҕԦ�O�{͛Y矺h5-d�ъ�gv���oA𡙞R�e��}#~ݹ��yg��Gvq~�ߡ��8O�{�\�+�j+�}G�5g��]��x�M�#Gh5C�Od{楘��u.4Z׍�*S�XG;��� ���$��^�	�m�6>o���8]��Y=8\����K&]^��:�</􀛢H�z��]�'2A�fȢa|� %�f�f4m�74V:��M��@9
u���g�m%�	�ԛ���έ ��J�z�`0�I#{>'��zi�2S���p6���	�bء��.���-'��V�djH�s�|f���ȋ\��F��bi�Ǵ���Td������풬ϸ����v��B�jc�Ȇ\�K�S&����jH'�������ʇh��A�wA� g[>���N�a���'��8��&qZ�