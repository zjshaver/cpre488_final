XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����S��!y��L�����Pnl�(<Vf;^S�|qjl�����.'��!�F�v��.�H�\��^��IqF�50W��89~�� j��ҢB��{��@������_e�47��O�#�Sf��q���J�[Z�(ٰ{RU�čwY��8�E#��M��sT$���e�Ô8"�$(lXgU6�{�Wu�OA���$��JWS�WF�h��;r� ���G���b��u�A��dvkX����%�},���@�yw�S��xD�:�-�H:��� ��	�e��ц� �!�h�{ڲK��?6gqP�^_�E�e1d�:GOL�eoVa�`�6V��>ͩ�6�w���{�Tt�x+#�A��[:i�6u.��ٞo�⨋���j�q����k�X�����G���C�������&�Vj����Y�Si��\����e׊�Z}KG�I�����.duR�Ek�`�A=��C�_���{���V�קz�.�,A���V����!�ÀD�)B�R��BT�}���'�|�֘�Q/�1FF��/zyp�b7n��n�iCԜb �e��2).���w�>�_r�����[e��w����ı�KJ�t�����?��5��o�˅���|l9t�qm/�U� @Pa�:��v��\�ې�`��th��!F��V�tD��}N��fC�&JL���z���@�9}�Uq���b�.���\�������� �I\�җ�$�נ(�ƿK�:'rL�ϓ�XlxVHYEB    1448     800�Dql�K��N
rL2�U�o��+T{	�4B�!W[s��b���qB���P٢r���ꐌgy9��p��S��&��L�VZ
���Y��Mv�k(���Y��6Y�v�L�T8�4u��\�
�C� 8r�����j���(X-l �cW~��X{} �Z_�XπU�C��@�vQM��G���p����������[hW����Q�W�M�^�N�ݾ�G��r��Y�<��v�S���5H��j�֑��AN��n�4�*f�� ������d�U�3�$�_����;��J��'ᕚvU���I��^U�Ψ��+�j�����r�۱�3��y�����{zy���-��-�#!_i�!����������H��t��C���/D�+fT[02�N�3ǿ��T�"P�qG���G���2/a�xV��o"���ӓ�(�&�8@ L��ז����w��zy����w�,k�5>�j��SE�҃K�� ��G
�4+�#�#��� �Ц���X�נ�理|nڮa'��'.� ��e���I�9�h #i�o+�g��=�$�8{�q��,jd������`�/�P: 2{�[��N1:i�����s#�y�޿W`[;`k��̴��S቏�E�:�9-s����k�3h�&����X�ѭ�>�y��I5�9��^;�x���2F��NZg`f��3:k1�0�K�fq������q��
���ݏ��(��N�X��>�|o��L�+W�+S
��kv���������"�x4/�:w���ǋ��d"1�x�]q7��W�~��C|z(������(���i�ȋ8��P_�V�Gy�=M]nLpn�y�~n�j�n��m�Nl��e�m������U�ƒ�j����!�<��Ab���9�a�V���bW`�\_���u%�nj�*�����%7�<=t��z���'��?�%�̛/�h8	�s��v��j��J  F����>D*����
�����Iύ_K�+Hl��~�B<��:��O �%�҃-T9����q=�_�3�Cy��-�uV��w�������$k� ��Ӣzy�����x~{z��4��	�!�"89Pm?͔�����k��f!i{Y�n4�Sv}�l f��gͰ`�j7"���t��l.��G9Lg�;������[A�ud
��5vâS'õo��VT�mԼ@f\!F
]�����As��Y����%�繐l超ERP~�_z���������@,U"[M;��@:/�| �v衑[7O��!�l�������-���;@z�Cr���bC,RW"=���SD)�K±,�U�2d���_���.ڂCb���׽k�'1��Ē?�Z�C0�����pY�PZ8��Ұ'�wF�@���G�t���)��e�ЃN������)�8t91�����K"�l��z�z���MCr}����b��}���ԹK�)�3A��^�ΤX�r~��j�D�h��N����
'w�i�zA�,]nz�(f�xA$���� O���d���6�\�CJ{�M�W.�HI4w�ji�=D��"�TE�?^����n��3�UQ�����+����/��}Ш�7��׮���dyZd��l��#R�S����l�� � �3�ÊE�z������F����3ݭ[����:٤���F�**g��lP�u�C7�Zn�.�+��d����4(�*(�&�s5���d�	�G�����ed3���f�vpL f�֭�7�=�׈�x�<΢"4� � rl�����P64�H�$�̊�~�_p��0j��M)d�V.ںg��o�8R�I�}5?O�7PP�:Ob�yk����Gw&I���f/���x�k�J��C���ܙ��㿡Cy�����?;��E�����BV�
l�0(p�v�SV`�@"�' �4N�n��?.��4–�&)h�r�����4x���R�����t-���#�5��θ� J%���y������hN�.��v)UG��-�