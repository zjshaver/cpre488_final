XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������~t�Y��-��*n�����uۄ�f#L8�-;F#�&�h�S��zP*D�����n 5L,���	��s���)t����:g��>��oc�T�vnZS4F�x���l��6IU
	<㈔�C��EBo#���`�!�����h�%5aDV�SK��_EԐK�Z�e,ʌ|Ǣ��o�.�ۙ�OG�J��o����#��㓞�r{Z���'tpr	t�E��u���"�������Pp#�3C������t#���nF�Kw�>؎{�� F���������̏�|�IDO\����CD�G��ID࿾Ԧ�|8r�0sd��
����ÿ���o��?�<8sme ��rV|�h����g�+�XE�H&�m��&�J*�Ű=�����5m�_m3�	M�Q���E��b�FK��X%Q�����[ȷ���*�t������Q����^J�>뎾;�B����Z
�d>����j�; ����?��}�#z%����t����#=&��F���t��u�OH��Ć�x$��"tJ`�M��n�@�d�!!�h�jZ���+�^��g�H�c������Q���ƥXS��J �uh��H�M�E�y':dB��G��x��Ldh|cP8�]���]*�ks��T��9�� ��B"jk+	{w�ܙ��ŝ�EY�B<�f��ESz�2�h�NVpke��X6w�(R��nM�#l�=nyѬ6O��cĈe�U2�\e�Hm���s���钄�~dXlxVHYEB    290e     af0}ST��o�/�~=�e�w1n�P�����W�"��s��A��k{4A�Y�|�ߔ��Uk�Ι���7�{af�C��7`�mz�����4an zV��)��ӄ�:ğՑlh��8��ՈO�Gi��=�SL�0H����$���5yĜ
����Amm;`�1�c@���#�&4h���6	�TEG���ƭ����V��s�GQ��Rb������톍P�G����I��apI �UG
��pP��O pu��iˉ�b�^b�N�ɼkVN�6�롚�$�?>\)j#K�y����w0�`�,1������E�#��ezp�#�|8�93����W�b�X�����=F'yq{��ʏ�����;��rH$ɫ����p$"]�,n������b9.n�F�O�}�6�&��40Pϼ�=0pFmY�{]���z܆-^.���[-�E�c5s ���6Ȅ9��(o�G�i߄:� �3ә�@U9�,m� e|��u\@�Վ�O�t�m�f.zL?!�Rgk�lN����mi��[k�����|�ru���5zu�ԩL�����t�jblt��������%5��i�a+�M'���J9��ǲ�į�4:��C�t1gv����!������T�QA�����1�'1*�;��"Y������;�9��E����́9��Y��<q�h]O�Wc�Bq��\�+5�,7]�%��'���MpH�"P��Ƕ!��O�*/���|��d���\bQ���r�~�Q�ȵ�ٶ�"v+ҊѾդ�������x鰹dJ�R�$�#� ����Jm�z���Q"}�-f`�e	�{,��l�a(��~�>����:sO12��]��RV��R2�F!��I���0iWxU2��@�!���'q�H��}�k�7t5�R�^5i/4��z
�m��giE�,ި���W^� 姢e�x��AiF�`�
�ʮ����F@�n2����8X�%�}𱴯����hwC�q.'���|0�����2<w��Dh��9��v{^=� �O�J<�S���W0EE��#\�"��4�6�|K(�� #�>Nɶ�����D̬��Dx�MI8 ��d�}�jBm%z},�/晛i�����Щ\x�\�j�6�7���)����(�v�3��!�v��W�2��zT���L��t��
��������������w��eH����e^�zGh,yL�.|z΅HJcu�<��>���b
e�EЎ�W1�{ mǩY�߬��2䱂����)��a[hkI�EF�s0o��Pі2ct	Z���^��GjK�r��e2BD�hr�;`eO�(Va�ږ��2��z� �-�[B��RBS�4HVII�U��>��bx���9av���{��"��j���;�q?�p,ld}=��.��臠`����g�H�ii�p��a(�W��**qx�M\��]�a��+0�3,�'T�^�uC�n��-s�(>����ݳ���]����d�L�5���Rw������[�wz�����.\'J�����CmD�s\��B;���f�&�x)��h [�}�����YYhw]����N��95Q��^ɀ_8���JplM�6#��P���Dv��K���.���6��ɖ�Q�5K������}⊳~��KT���f�E^=P��qݰm>ⷪ\��4�>b ��F�R�~Ҳ7c���;�_��#�fH [/1W/	2;d�<�cߡ�&���`�.7)P�s\Snǒ����}NH�u��\�:��j�T�&�㒭�`�Q���j���bG�!^�'o�*�ZUO6[oIR�GNP��/=.�F��%RK�t��xz��O�Y�z�s�@��d_��t��Ġ���u�Ӽ��]�)�bMU�b6��$+��N-&M��*���?��lX\�#Â*�E:ޠ��<��Fgߵ�J�~r������ݥ���<��̋�o��/��XS�ϲX����[�*@�%�=B-�����y(t�-��_�3������0��D?�uRj���1�NAڍ�5�h�����7�@�vEH����w+�H�ЋAG�*?��g�^��Y˖�����FBe��C����U
��@�P������"�drT�X�/c���-fC�u�S�����`����Ò��?�XL*X��ᙼ�4i��z��z����1�C~�݉�ѲjfT���_q���(�X7Z��`4�����Q��Iõ6��|� ��N��a�2�p�a󐬻�=i �p��k`�C	έQ!&�-�&Y%	�X�jO]�|�b�Dm���r::?.9��Ȣ.�x���� �HiZ�  WM��x�Hɠ^�G�SS� �((=��J}L<⢓���.Ǆa���#�}fh��*塹]0�{y(�ś�tC��#H�䂩��n�0����ōD�3Uޟ���?ₓ�����B>J�h��x
��V4�u�
��3��k����BA#zaJ��iT�,�#����x���ث=e6��3	%�ҳ��-eȃ���%�#�vyޟzmq!r��}����l$~�����`�ܳY�zrxH�EJ�ڱ���6g�c1�@/����_?��1��ic$�7U��p���HG�6	����Zy�,F&t��<j���	�Bx�7�n�)_hIһ�C�Ќ��}ٍ�Q���X=/�(I� ީ՝��2~�v�������es9�D���⭕;�m;���P3��V�L��%
m��� �pZ���h