XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���a�%r�^Pu)��UwzB�x�yƔPX��R_��w?�0=HuϷIv�&=| y!�M�m|���O^Ht�31�efj?��@/R��N��.Az�����j��r�O�7�����!���T}�iG��C�pp���~����ه���?���?�0�7d	��Z� AU y��5����O2�#��
�)M��8�MVy;��U��w�{k!��C�����oGB�Z���`T�3}j3cs������ߠ@���f��}7/ �?���%)u�#xb�j	���i�M-$�38�
�<��.��_�xS�{>E�&oDz3�M4�}�D�=ǂ�V�xP�����A�.�v�L���>�O!�����׼��Mv7���h�.�чi���+c��f@y��� M�P&���HA�� z�;#�x9�Bœ˟�n*q̓�Kh1�#A�m����h��d�)�[\�!:à�U��0o u�wE=�6B$�r�3�\m�ԞZ|t�yYFS�U�6U���Q���?quǹr\�d�
�]�
�i��{�*�)�t���v�iQΐ���)�q-��w'��6�8c��w���!��I��iu�����#��T'<��KM�p�Z��I;�T�
ey-P�Ȩ�-%g.�N_��˝���1�Ka� 6I�AU�M�m����5�ޑ�v�x�F�r��ue�=��������E���X����e!4�o�
���ˡ�U�P.B�ESA`�����(�eΛOB�Y�O��Hh����������XlxVHYEB    2b75     cd0���s��F�ĺ�ϸ�E��ܯ������� GXR���?O�4�iF���y���*<�?x�ɭ�
��[�$(dbBsfx�R~}T�pNu�Ӳ��s_�e�Y�Υ�e�������-C<�W�2at�*x	MJ��-��T�P��w���^_�2��
����a\�~�<�����e�X��[w��;Q�\B�m�	=�;���%Z�(Tխj��W�Ɉ0���[*b��(����b�Т{Sƅ���\����߶��= �>��#8��
����	��uZ�.<+x�?S(�k���9�%�'.FD��#�D��,nF�Aͮ��|����L��T�u�>|p�b��d�Iz�6u��ڃ��m�ozL|~�&kC8�'jc� �<���%�?WN�s����7�;n�6�&��#A$�� l�S�<AqBǣ/�;������%�Ao�ʡ�x��!���&��O]3�)ur����47$�43X1"�cx�J8��d䆆�˜A+3en�g�������:D�J�-�US^����9|�
� �{!UYí��QexZ���l3�c����h�&lX"[�o*'V����p_g�Y򚝛~�
h߇6E��%KE����O���2M�Ajʒ����s�B����i���3�3�(bt���b��(�*�֠o����ֻ�"������ڛC��B)�V��Y?ꏦy��}�W��o)�'�Ǜ�n.<.7i�!�V3�$9�c��v���`����ȍN)E5=�<��ǎ��[V@uT�_*~�Y��Ź_��q����W��O�%�q�P����B�7B���(W��s�qEq�j��+�L���׃^�����ר2�4�O6	�jK��s�&辄�G��B��
���N�c /���	�I���5l9�B�X�8ě�4N�t��m{.�u�a��'��A�҄�n=�+1�
I�R� �Mrp���Y�K�?}��B7GO�:_hHGk�h�G����6�
� 2EFҾ1�Z+�T(�/�/�t��WG`��",O^	��g˦��.����E�A�5vU&��S���C�R�j��I�h@h���w�	����xX�2u�{u�mH��̨9�w�t}���摢B�
���W`i4SM�1���/K�fr�t2��~���5����4����;6��P- &����ԹP�],���2��\ҙ�������sb��.����.ֶ� ~�W�U?j]��v>7ǈM�V����Q�H)@�2�LQ};�%����\�ځ��.6Bq�˹�9�����~dXj�V�=�-%JR�$A�BKm7��Ew�>g_}(6!ws&pM�uI�W,� �m�]�6���e9�@,��R[���H�� ��(�K�q���+}�*��(6�����8�}>���!a��QDv1{g���1Wuf�����
��t��}՛]��]��uG�rlu���>����O�ߴ.�M'2�e�&��<�gu�[�:�C����h�|��4�?��#݌��%y��\�yx���k1����Ϭ�O���i�����>���e��6޾=�>*h~\��D<�4�)��� ��d��R�/���&������Vm�͉��i��t��j��롴@ �@,1�k�U�S�ϊY�y�/�A�O,�1u�g�n�ӑƸGI��)o�Jֹzև�`�Ѯ�cx0�����hW��u6�k���j%,B�T��=�Z��7 �A_!�ఆ� L��@F��",�� �[�n�' zdP{�s�b�GYEОѼ���n�G��(�4��-^�^�D�{ʹ�_[B������壙3h�ބe��ߦ/����(,���,1*�ܰP��,�	~���1N1���&��:1]���h2=��ќ](��Kk��RvW��!(�y֩��_�s
�K��TL̘S	K�w�Y��23���k���a5&�/ �����{�%�FzUӅ,��wz�?�O=����Q7���/8Ǐ�,E,'N;���}���[i��m��c�L�֏ؒ�z�A� ���  䶈T��.;�0�����`-�wQ���IXa��u̓8滛hA��|�Ʉm F ��U1Yq��P3��K������*��:�b-;�K�t���h!��߰�(��љ��*� K���PF���*["I�i���v�Y \��s+��mtn����#�!�U��Y?���ʾz����d|`+3:|{_twP����z$�]��Q���V��VƘϸ��[CtA��_X����#=�}rt�0�-J�B��;(_M�McעS[�l��dT�)#z��6��R�ƀ�pM�Ţ�Ų�?F$�r��m�����������5�Vd�Jمh��*�T`��EPg6��S�,Y6�I�vס�2.��{�z�:BS��(�k�&�18����Y$���Z�@���@�}�V_Po4I��>z�%T�QE�E��R)��*�J@8��(�zQ��k��e�w�������������)n�����ˀ�V�PeHES��L�����鮊���w�ɍ���y���V�>!�����f�%�c�,u
��I�P����V��=]	˶�(�^��P�k"�,����b���DF�s�?.��7�"�9Ab�	lU+���`�CƤ��1�Ai"l Xe1J����=�#�.��H����G�4�(����G�҈f>���f�\3}@�$��/R�<:�ܲ��*�@�!9y��}b��<��= rvS�T|Wh�����69�f�/:�6��Cak���yw���O.L���};��2�X�K��4p&���<������b�]�S��jl�}3� eOn�;�LL'_w�f55�[�&����Q�xiv�����'Fa��#�ؐ���e��>.�2��g�u���Ή����X3�I�����'�
TUâ���t>\���ϯ�]�C��2ȩ�N��D>dti�|u`���V�ڧG����7��g��W	�QҶbt�r�e�����)�F�ĵg����L�B�� �|��: :Է�e`�6�*�+��zz�l�.�����)��KB
@�x�w�4g�D�������a��sĜWt�p��]�� r��O��ySu�Z�K�a�7��_IܪBB��(4���X��bun;lQN�#������$Iw��\ ��V9m>��SEf�� �CY:5Lr�X�0��^J��.Q4