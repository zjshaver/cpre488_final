XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������5b-����ޏ_!�(�~�<�
]M@��� ��F9�;�����T*�o���ٺ��q�O���+�t���By~��+�yD@t���;`<n�ģ���<��;C�`:��(��3RGI�2 n'�xe"jX<��W�$�0�G���	�������M��:r�I�К֧&r����Ú�t�o�/���]����}!���2�s�:�A[��e�����N�����O�7�X�_h�U?
�b3�(�;Y�X4�z�}�V�yíZ��tN��fi��f�n���z ���aG��S'�)�S|�%�O�����'�*� Ib��e��d�a��ت�����;����:��?W ǓȬ���"_X ?�m��-ҭ��8�!\p��u��ʚ�S�ih�"����aN��I	S�/��$�{��=++Nem�z���S'��LR\4t�N��/V�70G���ܞk��C���e�V�a��&����K����N	c�$h���\���i����,mb5�ܹ��尴s�&�L�����E������.�u�\&�������N��_g��b�?�u�7=�	�ǌ��?�l#�J��"��kf�~�ᨏML�ď���<�{�ޙf;9�DyF����۩�P�������g������ĥC��3��E���⨞"39�ݑV�����`O���F��B�;`W!�C"W�"z�&�F�X ��R�0p��5w�ĺ���2�^��3@C^`/Ĉ�XlxVHYEB    fa00    2a40W�x�z��^�qb���Zd�O�LSsV��5�D�Zݪ|��x����`h�oI�Y5�y��.�9����|)Aj�q�ĸ6�Q��9��=X>�ڍ���}�F��)���U����Y*���r��P�A���%�Ъ���@����9��4���<��5oq!�H�ԋqN`��6�h��a����.+��0�jl��:]"�T�y�_��uB��z��� ϵ{ᆀz�"%�t������MǊ��t�_Y�	��f
g^�a[�t���ӜU�rnVCY�s5ߠ�# ��
�u����q����|:r���<�W�����%r1#*�F�Y��7_{� ,:b���Lʊ<â�N�"C��u��UЫ �`����`/�}6\�gM���ψ��*!����G���vY��	�+�w�+��b~��йC�@}��u�<3��=69 ^˂�T��iN�>d�=�P䑣��\)i#}YF�'��s�m����	C���_�a�`��VN��}���p�U�7Sy|Q��#��#��µy��^��ź8Z)�`f�l����Gur&�>�sU~I�i��{�+�ȅ�:#R
���u(�H��� I�7o<�S#2.�nm��� [���&Ve����D���ȕ5���Gt!�C{���E+�<���P����k.#�^n;��@M�B��R��V>p�1T�'�<O�$�8��mtg����� �3ǅ���=�"�d�>�˔E�1��B]�d�;���_�i��51E]����Z�u�`Q&X�K���og7P���LSL�j����e��9R=���J��D��k�a{�e%\$�Bp�PuL>�O-�����٠��/�Z�J���ܾKKJ�ᡌ�eI�c�����f��uynec��J�ل�"�م��\�"1�-��w���8`�1�}hi\#��Z �H����x.���8�؎�A��;���^�$�4���R�rlg�E�Xأ�T���e�j�8�G�O��
��dJ�.�m]�D�����뜮P�1";�y���̗��1Jl$���c[���^�j~f�Ӓ4����m�o��2�kbM���S^�nE�]~f�gp�Y��E�}�y��S�����Y
2��L3*��\�o��Χ��w�9��UL�~qa�9����ʻ7$�M�^����/bC��^��S��Xӳq��_��'=�5! ���]����Ǒi����������
~����D�F��}g׬��Bj3Z|i'tV^��9�%6��� 9Y���Raf�A3�ˁ�$x"=�B��m�ޜKB4�L�ܵ�n��ia����"��S�}V%8,��.g�/a��E�/����� 4�:.�S{����������fBF��/e���*��T?��O��}�����)L�,��̠v#��"�'}��i��ĉ:S�|�l�ί����àE���^)�������1������f�{�
*����p�Z}N>�1��z'����p��8O72��Z����ZI���tyRZY	M��V�f�;Bta�Z����8{j����X���q)1��*r���=�K;��A  ���${m|:�(n�3A�.U�T�38ri(�Ns"�h������finDAOP������d�.�y(x�o"K��+�#З�M���gMI
ͻ6m�_�(iob�f�w��{jf�^��˸C�����_>�c�\�gB��Xv
�
��q�n��3�E��.�G:?���5�����D\�I�ى��op���'�N`ܕR�d�t��,:''�F��.�$��O�'Vpc��c{��ʩ'�L$ď�ۉ���Ey�K��(Bn��?�����́��r|�g�?�0������{9O�8s���#���ĿͲ����aXix1�X�Y����#=p�A[����� rѹRd���*�k��Ĉ��>���9���5�0(�CQ'o`�mKI�u�?!,������ѝ����#s�ڍs���4�䯖�rZ5�W�w���q�XB����:�������{g����⹊a��#�.�S̗!���w�:P�9�Fr���^PR|Fc���K��J�*ĸ���؏p��A������TѰ-i�7�A|c;i��.�p��*��6!��o"�0�W�$���$N�'�+I:���S���Pi�+x{!�`v*̀��c$��h��8��M�7��%Z��_����Zg�3{s1�g�+P �������N��1"�]���%1��2�彨ap��4��1Rw����E���k�9�f��&���a�[�:ZE�����~���uOr�A��.pr�ަ�M�Nr:����w�3�_� �wƘ!���Ґ��ޅ ��U�p��4�7�
Wo1�/'~D 7�C��kH9�MHr��1�V�s�߰�D)�ARg��)Cz_)K��V�Ȳ�Rl�R�~�KO�<��\�]g-:���LN1_jzMv�W���O(�_�$��L��ގHzB%�2G�R���xݿ�2po< o���q�����>׃|�ր��+-צAcM�0-����A&p���M��tj�����c(��#oUR-����u��l�sgm1_G�#�F��-+눲��R�~����O�z����ϓ'�C4��8�|��Cs���@#/��@_o^2Y<��z�@��҉G'��	h�<X�ⷒa�B�~i����_g���eZMJT�ǒ*��q��`�$j����嵍����7�+��V51������&BeF!��K|���a!������s� E�S*��5���'��R �!s�2��ϭ�~���&��4�?��%�֨)$)�ț��
��ٞ7ɴ��XS��_�.=��P�O�AȺ���3����-ɲ��ca�5y�Ha�͙X���i�P��w&�#���_�K�����鹦o! ��4�6w2��y����.�3���OiL�Sɜ��|<hz��=ȣ1ӛ[c�ņi1Ә	B^2�[W��8-���Jh��>�<��j�{�Kh��,o�N�u��Ʈ4�]��|W��YG1�Yޗ�ƥKF�NI���������2]�0���̘��fw1���
�
(_�*[ai�z)�6�� �!����'><d����9�x��1��{��!�i�d��w|�@��?��U��7�8�b�ɟڅ�1̚8c��zeBXaB�Tm���`���1�W��h��Ȏg��#-sTx���
�Q�L��+W@����Q���,��<�.�'��}���ƐUz�ݦ�g[wr��c�-�o@�DSk�	���sn%噓�H����c�E4���6n�Q�����W�䈧0��V$�jB�~����#�-����s��$��Qa$�/c�^	cW���1aihR+�2ǖ"Z��j��pDՉB������%u�.*?�^}���?�"3̺I��	��y�ׁ���k�j'Ѽz�(3�en�]X���t��&?�e���$35�����F.��H2e��?1K��e+~��/���ú]nb���,wbS�&@� �nAn�f���|�U���*W����Z{_��beVs�:�mL�.��޼f���VVDorݜ�T�y�?�7�8�Ի�_�U�<�'��c|�yG��I{( �-�t�orO�#�`l��ieB��ɍR7���}��'���R�T�3n3\R�1�T�~���*��!��f�\�P�a<^i��E�G�� 
n�f�6؋��9f;[�۵��m�]���ءw�M�NA�����ǻ��
������֝<�0����m��=��
8d�v�	&\uX��_�����j2a�#1���L��*Y_��rx����9��k;h��o�I�'P�)�UZ)�;�({��Y�W�+f3�����H	^�y�s�gU���'0��H9p�W�<A�a=��

A�5�0�-擥�τ�s�&s���Y���g�|����N�
TT�_�u�}��gH���.TWLE(�g�������-��Q5|_�!F�,��ͫ�����$v(��6 �^��E-[�^���J�|{��g��M��=��D#�ؐ����B�|��A3ɏ[���g��D�5s͞��l`ۙvk�l�Vޯ:~�M%���Z�Z�@h(~�U| ����m�RXp9�B�l�^D�.�ˀ�Ln>,"�y0���x�l6w��cU$��ϲ�� 4��CR8����H�yug8�����:J��8o��)��v�����6Z�r�6�b��[?��ة����`$o&Hƣi4d�3M8��>�U������@���KmW��ˮ#&.O�a�H|I�:�E �g�����1��� S���ZD,�	�ȍlA���/��b�{h��sf?��'Q�T�?�wd�Ej���ߦM�vD"Ơp�$����>�r�7�WE���t�$�0�5��ʊ)W��-j��b`��v��\7�Gؕ$�ѧ,p\y��ٰ ]~߻������T!T1�^a<�R��h\4�����6`#�~���Q�P��2��?y�����ukK7�
d��V
�'�S�߸�[��%�\��( 7���XnWI��ǽ�i����j��n~��`O�Q�I��ܔ�ON4�䀬�y'��D����ڭ�اy�C�/�9%�U�kC)��w8���_v�)-�N?�Ƹ��_6��Iz8/G����f.�p�`��~ox�|���u��0�ʛ����\�,�Y}m���V$�t�WZ<�iWR����{ݵ�Ͷ\J\5Z{��U�C�i��ƞ��)�3��ɭ��C�U�%�۸>cpw������L�M�'R6ldUh3�#�ԛDP|�o�e��i���<�ӣ���L�Fũr���y����P
w�
��)�9^�U��?5ג}||���f�G�8eV��;$lu^���.�aMJ��rB��g��?2MO��R�������"�s�RN�rH��jb��RaW��g�и~hk�����p���� �J|
�N����_,����|�rډ�����{ѻ�W<�=��y8'����p�GX#� �f� :pXWI�ҵ��{)����r��� @j[��iG��E&× ϗ?5~���rߘ��`HĹnY�7Y�,�'��*+�÷<6��ƅ~#10��y��M��U�}:��t=tIŰO���!�[ܱ+n^Q?���|LU!�ɾ�;(E���ٰ�|�)��\]<�i�x�ͨ�x���%$s�@�إ.�;�g`:G�F��^�ȟ ��VD�Es#�j�Y��7�=H��-kQ-�s
��P"�4	?�d��eV6��e�?�Ԅ�_d�����E�de57�z���sb�1�y�k���`�{;�����<�P���'1�]�(��-��n]�y.���8s����.��tv�A����+���b�Y~ěl�r���q�ҽ�x��z����"�A&)�HX�(#ed'���B0jP�$w����	�ѥ�$��5�1+�_�V�/�N=��-��E,�6�I&�Y�U�ۢ��h=��s�W��oj�p���_txԍ�1��cJ�L�T!c7.��U����`ߌ�����*Z�ֈƘ
����@[c � �vu���	����>�Ė�&[e8H}sJ��O���;�"��.>AW�	�����t�B�%L����NAe�?]���H]X��W_��+��.3+Cq��lDc��u��ˎ�g����i��a��#v]�EX�])�  �F�JdM���ebw���#�f)��.�<�ܨ�(*!��b���7Y�A�����c{bO��,QTq����p����H����ǑD�ƌQ�h`�O]*�K˦摁����|KRTH��0)�,��9�X�u�!J�߁C7C/-(��"��i�z��F�,)��(���MQ��Q�(=�+�����CN��`_�M� }��nQw$6@�������jؠ_�Щ�*$�m�Z��E�D R+�=�ԇ�N�^�c�+ҍ���΢A�(��CS�A�sGtD��dS�P|Oq��F����W2��x�8��V�J){#G�ej�du7��0�
Azk�v��Į�o�мp0�kG4R�ڎ-��`��x��!� L��f.�m�N�s�U��=�2巅�2w��\�|��t:�����0s�bY�nW��0�, y�_@�&S ����o��K�#�M����m�	��&&�����\�'���9V؍n��vu�7�D��d�8�A��HcHf�dxM���m�����a�\	�<�|�JK:oW�J���\���6��<'U�`��ZE��\�J�5�,���,�ޡ��Йf��p�At���d�9���ցk��_(v�� ��� ��s�a?@�2� �ʲo�V�1G���Ƞ�@D�-����ڏF=�Z"�gE/�E?&��Ԅl��wY���^�@ �}G�%�$�v��t�c0���35)�Fxuc��q��?s@��,#�#7rBA)B;�jD�CQ<"��9�c�W��5D3��"�4�{��;��� �X����7⑳�����ss��^�4F,��߹�#�X�ܣ�|�R߼u�F]:&��S�mh���Y�q�O��u
����(֣6�W���W���Nc�	 /�����)��4��$:�9A�|_������MUE��7;m�k���Uz�q����J.��W2 �,_���!,���o9�[��M��������������;�ɬn��Ef/
���>.�]�o���w�z�*z��e_��-s�I ��ޔ
��]���?*b���TF[�#ݠ>u\p�J���~���ay��f	c���B���Pj�m	�����Es]W<�%��D�x�m-�f?w��S��y;90�^R�	<���?j&���4�3:^L�P��I����U��2�@�
tİ}���Z4�-����a�z���5�Y���Zr�T`,��	�b��Ch�}m%�P0��DՐ�Z��Dq`ʳtcE�����#lb�r�,�폅�f�=>{rԼ=��Il���ܪ���P�.(�F���!V��� 0nz.���lZ��V{�~�~i o�i�2f6n��\�I��8܅�B�u������8�75�nj�Х��)��Hed�O�TYV��.�6/BB^
�����G1Sf��VA����z��űun&\V}T.��X�RN1ͥob�h�J;�7�^�T;���ya"4	Ģ:�DY�mVQp5$p��9@�+����&L1�f�Bɸ4N�Wr�r���f��#�nZG{LT���m�vi0.Ts���ej��z��K59��ǃw�t�ҾNz��&dD�߄) �*�9�2t�� A�xڙ��N,�!�0;�Ԕ^��z��~�D�c���I44oJ��袊�<��E�N	,O�D�����R�M�/G�[�|�(�~JgHߓ5%���HSLQ�s�g�î}�4�f���lS��g��N6y��S����y���rao�>:V��ǲ��� ��9�ڻANA�&i_���<���uq�ӂ��Eb]&�� xU{g�6n,(%�dW�|���L�����NE9knF Ə�����GZv(o��7�^_.fz�:��]�Q&+'��΢w+�ii{1�#�s��"� ��<A6���	��{j��H�s����`(}����Pl���_�X#���p�{��6�i%��n�[��{��fqb��5���4����moh����o��F�W�ԮZ��Ǆ?֏n�#]9���Q��U������2$�uר%!��I�S[�P��~,5볖�Z��i���7nF|V昛U'��27��\<����'�j�<��"^�j^l�2�}N��xU���&�p��kfPi��K�M�0r#� ^��۴��f�=�pU�I�uS�4ؓ�B@�!�Lȧ�� 2E�ۤ����r�_�J����M��Z���XО�9�m	f���5Y��"��Ykiݒ��,���ϙ�OӖ"�o{�L��62�W��0�xݦ´d�ޓ��2��G~q�Ȳ�4�Yܯh�_�}*��|ķ�YP,���a�a����+�������I4��U}��f0J��GE��Q�ELr�&2��P7����#g[C�d#�Y�JN-ȯ#����m'8i�3�ْ�A[�/�`���Oowo�'�c� �����'�&.0��$r/?�#���[��E�����/�N�����/7(��Xr����
�ܩ*��D5�t��J���:&	����q	v!��{#ք7_6��By�|Y�.m;#ަώ[� �M��K�;$?�e(3MP�S�o�.�8Z ă��;�qs��$�V0�o������*E��z�m�zN�~��L�����M��~oW�L�~�+��F��Ff̫Q8��;���\u ��]��ǧ1D���
Ԋ=E-Ź��
�2�gF�l]ס��QՖ�8�ޘyɵ�>1r+C���ꀨ�x�gt���������
��t)","lF�R��o�pHe�/fE���=uDsB�?�3y�l��5r�s����$)�g��V��9�/6�j3������B-	�E<OC��p*3��}�9g��xMz�̇fT֌����?�+k�NWb���/�ח�����ӣ>lF�=���'���'.3WN�O'\�V�>��*f�����t���i��M���}���7�����6I� ��Rq�HO�ݎ�b�<1%d|�����V%)��./y
fc�(paB�	�K�6��I'�dT?�����y�G�k{J�������.�Euv����[q�.h3
��Mk6�P��PX�(��E��LQ"ϐ%�h�#�I�	�W��q:���[A+Ǻ@:���B>�I���wDj�H�x�U�j^{�Fǫ���nŨ�p�͟����Y���>Y0$�4��ر�!J�T�z��E����HT�ZY�5�G(DLYH�P��]�Ke:�mbh֧m�)�yǷ߁C��)����=,-En�u�f>��I��|��!�ʓ_�ϟh3ezM2�9���I��<4���±M�uK1���5ܼ�t���%�,�;x�/�-}b�wv_{�"�I7��Y`b��7�Ɠ�.0n?����)%�1����M�5��c)A�DL�x��tu=���Gou`�������i^02�.��1�9�ǂ���g���B��%���3�Q�u$��e�'��L�� ������z��7u�jZ�ݵp�V��$�n%c���Ʉ	^1���ꃈ
��[%Gu��o���AM��T�Z0q��Ո����y����Lh;(��6+���*ˬ%hN}�#�ֱ�vu�{��[!}�ƪ<��°H���6+�oإa���oR��<��K�-�}��l����E�Ƌ�M�� �gU�hE�}l�	^dYY�����	"+k���������)ԇ(��-�8�c����n�R����E�^ߵ�/e��FϴgP������r�m�����*��w8���ħ�ʱh�^-*(J����K��D��n�)�AC=�����V}���2�< ��J��,�)r�S8�6��E�1B��&f�O�*�C�ҷ�A�hC'BA5�O\2��~�'eJ�c����Y���D�A=
2����Oसe�z��r��7P1I@*�H=���n[ε�lT/|Ĩ .��&w��	��9�]3�'M� 9������0vda6Du��j>\>U���_�X����W��Ru�V�>Q��.����ЁGzN���A�+��7�n+��с���
ځAz������/j���������m�|�8�~� ���`��Ϗ#F�F;�^���6vيO�C.���[�0�=�k49q�����b�R�����^r$O�\���M�A��d�#rj��T��0�J���?�9� d](ʼ
�8�T ]�B؄�ևh�yv���K,�Ȣd��8o�\Vk���nަ���[��0��g��"W��4��0?tw���a��?�֛���t��ɽ`Nu2�0� )���sz�h�ǳ��S��{l���_�T�٣OU|��ͧX�k\�e��PQ#]�4KO��B��\����]Q���&����d��we�=^Y$�������_Nn�����f�Q.B)aks�z�4 D4�-^�^tL�`�%�[� �����2w����䏁�-H�a;��*,b�w�} e%�٣w�NAJQ06�Ƭf²�om7F6��t�d.�Q���-��lO�� B�=�wf�,ie�x���j6������n;n{4���B�i	G!��rT~9�����'i����ÑeH��	Ы��~�����X�Zl=٥셹 /`!ݤ�d��5h����x��o��v��c����b�EðQ��IJ��p�?��f%�3��auUx�=������K�9�%PP
��̑�DC��l9�0��.㛝�.}�煑�D�>��[���FJ\<�xWx0�Ѡ����J�Ȉ�@N��X�?1!L��	!"����?�F���E�t�����ǅ���!H��6J7���׈A�������f7�U]�����+�=��l������Ts�A�8(�O��4v�˩)�+n�5Mܟ�Fξ��\���>�hZ�hn�7]���I9�S>f�3y)๯�'��l�ɪZE�\)�H&��O�~W�ʾ��mY��=��z�=o%#	�"|ḤnjqE�+m����L
�-Y���XlxVHYEB    fa00     8e0T��uԝ:���������&�P�(ǈl��7�dS�h4E��09�r
��G���H4&�Z! ;�!�_��yVVYv:��Q���e��0���[	�TQ_"��o��V���<�r�Si'S�e���I8G��a���=��w=�K�H�\L�{�-ϏN�t�����6 f��Tv�b`��Ep��/7�}d/ʍ3��?��P�`�k�~K��C�HS%�:�٦�ka��4/�Q<�5Uܹ��O-��̎��RQ��=�����Hۛ��̜Rn8ǫ�u�b���4�O�U�ʅ�}D�m'+��� W���ڎ�lMzZ�E걇� ���[�Wmi�� �P�%g)]?�3�e;!��"��&3��:ts��hlh��T��,�D�r��coo�1E�0�h�'ܚ�8LΩ�?N�,�f�	K,Y����	���j'��P}݌ �]�$�$j�� פ��AQ�gN�o�K��>}���1���	$���Z*�ʳ�$��0��a(S� �h�샘�9CS�f�=V�}3ȸc����f���5|G�\Ty�$�q{!/�>��"�b�6r�4V8��eu�2���2-:}�V�t0�OY-ѐ=�C����E�TM���n���HF�����_1�
cw!r֏aXO�W��I`�;9�q̻�ʸ@/"�6�T!�	��x�������#�ؚ�t�3&c��M��_�
*���u��#9�}�:�y�zs��}2e��vg���ٿ>����E�=�׈%/fH�|��P����OS��-��`3��gw�7��^RJt�ǆmo�C(���2��*��[��J��w:�G�������O���M`�y� ^.8��<�͍��S�ƚ�2lI#�|��pdj2^�r,��@�Qvу͠s��3������:>���㙙E�P���p�-�������.B���D�*N�"��f� s�.s]-�Ny����d��3W����cMpٙD��-K�n�Xc�(d>���Km$N ���Bʚ��q6������p�X��*@�@�ԅ��?�XV:D�b5Pޝ��3�K�g��a�lP3V��_��\�����vù����)K�Dʀ�/E}����� ��µ�A�_{�E;E���|1�����h�h Ϝ$�t��i�"Wg�/~�|a�r�GŃR�Jf�U�;80�}��Ѝ���rp���тV/K��]�cKmYZ�1�'h�s]n~Nf/���� ���j�g�ͼ!o;Ε�݃�'y�@�C����<ȣy�{�_�ݼ����[�:��٢�ɻM>ѻ�3@���!H��)���V���N�����%�~�>CG������j�}�^r�DT|X�|���]ejy.Ss�vͱO�
���/G�Do�A�EU �u�I(I��T,:��(����ut�>-ߋ��VL�|'��0�h���D�|-��u�����Z�������c8gɼ̜�ӱ�]	��X��#@���S�����׀����a_-�n��D|3��O�U1��2!"���A�:ˢ@j3S#�en�*�,��upzR%C�U��8|�T�h���?r8p`��2g�2UE�O{0�8B��A�	B"�D{A-��b�%F)VW�����Ѳ�3��B� �{]Gq��d�m�]���Xvy��u��§F�٤��0?�T(:��$M L���y����E��@�_����}�{ �c����� �6�ϽA��Y�7nLH*��}AH�n-�9�ؐ�|f%j��q��2t��;�p��k�qt7ѡ�`VK�_������᪕yE�S�E��.+�}\�{�b+�ͱ~Ui���c��5᳈@�w;�(U���O��lz��t�'j\Dj��%���Op�$��R�\�):!0������7���K�DXJf����!J���̶���#w��M������	y
K�c	W��^����#?`!1��LU"&}z����fm���!q�ސ�g�_�]������ؖ�B��`�'/*�6������t�x���{�q�^��~qG+j��x�����։R_j�3m�?����PZ5�o��2�}���^NXT�w���qBiUX�xf�TbD��&���>�p�X�)�!MY�1�����ӟN~״����@*�Q`8�BU*�f\�s"��x~#
��6,�\Z��1J�I#w�wR*Ԓ#�N��8�]R[��ƭ�?�����KmB�_�?�.7hyXlxVHYEB    fa00    1110�����/���.{�M{b�^�~��p�H^���d��68WO�����2 �X7�\%p�oJ�4Z�0�%��]�/ҁ�V=��&wnl�&�_�����ɽ,�u�tVؑ$�LN��Y/M���zF曘V�W�(<��#K����9n&J� ��r��o�� [��iX��rNW�����r.�1�]i�����f*�_�~��嘸�ײ���TV�R�e5������F�nM�'�ٻ�|����l R{*��wx�ʓt]UZ���=Lȱ\�Vq4t�׽���|���L�,��d[��l���},�aG�$@Q�9Q �Ǔl/�������_�w��G�f�D�O��u ��>�2�[FFX�����AJ���;�ͺ���P#�ÖY��؃��~�e�^V�麟����>뱐����wܾ� W�Mt�x7��m��({�2̵�u c��~�	����y�s�?v�e�B���5��]RYI�/_��θ��2�iZ]dxsey���,�M%���@�6���_K��u���L��$3�!�����$4��H4��(�dq)���`w����X�X�a��e��{f�+17�0��3��0��P��������J3�ևWR��+�IQ��94�éy�J�إ��4�.isԽل*��h-m�`�}�{](p�y�"�j�j5.^F��E.V2j��	���ΏǦ%:��V���6V�%�J��y����J+���#����b����5[�)'��z�0�����17W�Yb[�$�P:�%/���~�۔��z��0tA�l>�&�tӐܔ�<E����J��Ն�xyCy(��p!5g6�`�Y�b	����b�q,y��7 ��i�E7�c�|������L�2��}ɪvj�
��z~D�Xx�RN��#��QG�*��J�VV���/K�ɬQ*������d&�N��W�K�k�w���5^�:=c��X �R{�I��~[��]|b4B���g��;�λ�(�Hp�������B���Q�7�JI�n2���[�K-Vܷ=.���I팛Tx�u�'/�B|2V�`������Ȉ���%H}�}!�����Ek	r�i�B�_����1Z_��߸��̐�!���Y�D$�(4T�K�gE�& ������t\�=��'8�*��e������fz��IqMj\�c���s�@���R�W������AƔ����f�9����Х_���in���& ��/Zi���/�Y:�0��^�e
=ҊP�3E�Aޕ����b���2/��^!k�q[n9 ZL{sx�	[�)x��y(�*R���?lt?	�YP�����K!��
N�,ٔ 0R]��#��UG���/돷�u
|�CIng�������*9o�&��Y.����߮�	B�r[
�<h��]iZ=;Խe��#G"�)6�ы���B1p����U$�Eǒ��� oy9I�j<©CUh�=�`P~���s����<�L�4Ǿ��v:Χq�uZ�ee����Ϩ1���֦LE��+��dg3?�;&O'Y��go���u��[Lh����PU�?�!k�(��h��#$>�gd�P�ʴ�u�qǡ�4��A�d��m�K0�9H�?(����������z��I�Q!�����Kl�/�
�`�M��U��A6����x���R�����hX.t�#Ċ�ږE̴����,�B��~J�:�Z�(F�[�J8���1�B�h���w�<Вc����w���v�N�r��h���|�jUk�_�KNԌvqx�ӑ��t�K
���NfP��I3Lw"��~�S�>��q0_��������!O�m�h^�܏�+�Z cx�&�K��R�'�*�E�˗�t�6ܰ㾝��)�7����9Qѩ�{�c*����d�WT�j�^)Q!�6Ʊ������r"�.W�!��#5 ��� 3�(:�yv.���f<M�M��af�h%Yش�"�4*����K��ֶh�v$�^1��'������м=1U�����j��Y,�=�'G�2�K�w.DV�u�^WԠLٶ���"V��� ;Ց�-�E�b�3�]����uiR�f�lN��ɵ��A�E{$��-m�����G٭��7O�~>c+��<V������m��f��̺֥yp*^�x=��,���i�K�b��v-U:��g+x;7i�=,���)�@Ҽ�05�efY<�k� 	�`��It����+m���l���Tj9��V��~��fȟМp)����[��u���z6=:��v+�3q�e9Zt�'���JX�AF	��?4Y��y�ԛ9f�#�huS�8;�r�$|��z��B΃��Ő2s��p��>���RpD8[ߋ�,WS�h�������m���q�o��*6f���ĸv�1N����{\"��Ns��G�SDu�瑅t��iυ[��ޫj�#��!��l7a�����|S�$U�m��ۺa��f�+�.�>9�.�?J���b��u���jnnT���B����������V6 ����c�k�� l�U|	���t��Z�����+�>����+��]��s^�*-�Qtf`�[%u�Ӄ��V߅6?V
��m{��8k3��>��V����ԩJ�.�ܺ;��U�;��y����z_��䤪�s�x^.�<>E|�y�8���,���!��nV;B�uk	��������)2pF{ȆX�a^e{Z����3isQJ�@V$l�4f�_8Oq�= 7�)�GhJ���$���ۥ6�	���(;�����i�����b]��5M�lď���g��j_�o9���˘T�+�ԗ��<ʒo�y��юS8��*5�XC���+�N�)�z�
�
{������q�R1�]��a�ow毷q�N]��Ľ&A�A�ni߽PգN-�g���������)3�h1`�n[���$P�I鲷ퟑj_��"L�*�F��[=�?Χ�O0Ә�-��m�)3o����;���~�F���w�l�՟��W��t&�?a|��'Le�+ ��$�b�Ӄ,�����Y:&xP��ݞ��& ��n�T6ٵ�?6�*b��)��r=p�D9p5�ś#-���
f+��X�{��jqʆ�)*1�H��l�1���\ṆA	���Y"���lc����&�u��B��.�rI�G�X���/ak�2"܇� �2<|�����ec˺Oe�Ϫ���������[�S�Rl5�T@�h�����ܝ�,�r-�G~om�.���c�Vg1$���;��� ���u��Y!��q�ܴ,�?�[)�o7��A����g}����k�/��2g��w�(��lXV%<L�i4k� �������M��/����\K	�xt�D��<z! EK�>�*�"I]w�mD�~�:�*�eKt���XX4���F�Ika.OmD����λ�s�>���5S�l����8)"5��U�I/ �7
8�Mz-�k{�Q��Lt�C�G�n_R(��4M����m.����'4���� ��/?�[�.�_��Ht7g��]��m�J2���V��@��D��<]�r��i�{����Y�7b�b�,c<<oh1��u�*c/i��Yi{������HIy�E�P9m�ƤGh�yƜ��*���q*jL�n���(�^l8��[A��Mr��<x��'M@
g�:F���K{Vp���6��������(����됣��N���5��1�����1茇*�Ÿ�,�{�t��]��V3��� ��'����K�`���:R�N G�L��F��3=�Hy���Q^�ȶ]q ����|�۷�x��3�k|d�:�ë�hF�0e�&�~0*YT��z���ܲ� :��+��L�ŗ>䬴i�w�C�ڍW/�b�PL��=�|��
�.��P)e�?��LU/H��Kdp��N�xq4%�ŕ�)�,JS ;���ކ�L�0��<y�ɗP����s�h
R��W��<�\��'� ��3oV���e��,��_�#~KۍH5�9\&�����գp[˖�Ӻٰ �h.1C=k��M��6~�(L��Ͱ)A�^	�ӈ)qr�EAҵ���B��&hg>݉g]��ap`������t}�}j����v�M�d��ϻh�!z�/�{���Z]�ZUx;�5��i~�}�U	/�o���hoJ�[kE�£(,*L�V����z������м����F�ʩ�	��0�LI݀�_�TvGL+b�>�Jq)>W/���}gcZɏrnx�~���-
��u�$�V��v��R��ErN�� ��%ќ\���C[K�P���X���a��hӵI�?�XlxVHYEB    fa00     ca0zے���`9�*�/]�&�^C��Ș�J�r��R��"�f���7kg����b���3d��M��Æ�^Y������7~f.�&>�Z<�����*6ñ-�������8@i�hb
;�5�t�v^>���zZQA��wo�7�ݴ�+"\����~�K̒���[��p{��_DMΆC�D 	8ވ`d�3`� �*�- 
�r<o�~����RU�8P�	a�� ��+k��\;���-���_�i�ߜ]�"�,-������WXɭ�5D��*Q��h���=2�~������ײ��us7�+xX�y5�d0BW�4���z�ly��6�|t�T&�7�U����+w����É���&~�,��D�WQ�Ⱥ����;������ZQ/,�O��[.c1�2�l�
Po�!Aњ<����.���	� UMv���j�����PJN�$5}��gMSՀF0 8�lI0&���"/�����/Y�|���?�q\APvO��.�m9�-+��>��R#�X/���!����ƏrKjwݒ��C�Y�"l^k�"�[p)��/����=�ll�ĵ�k��`�B�Y�Y��5P�� ����Q�t���D�|+��4{���/6<3%�)����N�n,s'���/�o�t<	�TUȔ���e>����^T�9���Fg�1c�~*��^�f2�
e��0o�xV���H�kC�Ջ�JX�ִ`K0'�Kyh���,T4q���O�76f�#%�ud)D�]�pK��C�?����V�n:�vb?�����iYw���+���"M1�\��7/
�=�`+�Zv�D�᪫��CΏ��j�ecu5�� �|�F����J��y��|	{'%HNY8�9�~�F��ꅝ%�0�hP���8�����8�B?���u��@jb v[2�ە|9��f���ܷct �1v��jK���u��o݃�yȷ\;/z�ҍ�j~n�ȿ`UԉDX�n��|��kc�E�[>��y΍��7��O��n���f��Y�Q�I#d�'*O�H�i�Z=^���Ԇ�Mo�����8-��x��@�jwki �D_�Z_����yc4�T����>�z��P����v�5�5^�
���k���]�iyw�ko��-$c��kY�0R�b�,�����)�z�1��l���ѓ��_;dy	$}f��S��Η $jή�vz��p?��+�ߣ���Q�K���]��&�6��U��Ii� �Teꄨ~� {e"luxf���ހ����M�?��y�S�S��ڍ+������q&�gV���nD���u�giT��8��+yZ�v�.l�L%I-n��O�����6fM9u2=� ��Dͼ���h�-��<O��@@��ȟJ�ȫ������:ȢB}�5J>oZ�0Mi#&��`�h�ƙkD�\ɔ�0�z���J��+e��pj�F��t��Ƕg.4Y�Z�\��T_�>�kQ�e��Ѓ�b��m�6���O�|��1�A�3��SF��S\;�YpqgR"�l�n�k:\�d1c���d���1�utmO��*n]*s��Y�ʆٴc��ow�*n�-��^9�㚺�]�.����@e%v`)x�~�Vn�/P8���jv�xÚYϳ�q]ؤVU��p�?�c�B}=���u�N/�. �l�T�g�)qFI�(�>��<;+�g ��F��ࣆ�c�a��[����ۓr[6�$	%�:��I�w!�ݫ�{���9j&� ����Fw�n�O��z�z����-�P�zy�E�;�&x  ��\9�@�S��r�����x�F@+Ѹ^1g O<劲��y��F;3��l�E-~2����6JNc�Կ:�j��P�2�%^��'0�M�2Ғ�ؼ��A��T�ګ�9�b=PզE���}-\�xrG��=�y�=Y�I8���=��F�!9+c�B<�4�ɿ͠F)K����ڭ��<��4�C�%���$�0Xxc[Z\�2���� ��C
FJ>����/�j�FZS�]s5̀�b ����ɏ{Hжi�3z�@���Ħm��N�6�o��g�*hK	=5'����h��O7<�rHP	-�3�Z�h�J��/?�2�̌��.&����p qR����*��R�0����.K�h(g)��b�w)��G�}=�%l�E<�����b2`ޏf�7��ȝ��NP��sx� 5I�<�(�*}9�7�R�QP�j2�n#NgF w!B`Jz�f���D�����c"�����e�}ՠ{�$/�Ц�����#�R6U�HC��(���s��EJ_c���ᗗ�E�T��V�Z�膲���S�
7@.Xt!��ᅌ��^	ܻ��wM���x"���r�!)~"n"`o��j�2BM��SK.N�A�J��Rl���� ?�|z�z1�����j@ȭ^ŌD�
�9�P���������L�`�&i+�H�RH(2�Άn�{�. ���ߝ�i@��>��<ץ	��J�z5q�?��ZyR��!!1���6�a����̩��%��@������*���E���K���	lz��̜־��wt!��L�|+��.�C(�ih��b&�ϢL��HE�t�Z$ʙ�$�m�]��?��Vn���W'G��g4��{�_�Ix�T�
{�U�P���P�*ѥ�&	?��nB��n���P�f}R� Ս�bS8(�[�r��#����v�D����m,>ݧ��J�xJ�sG5�)-��S��*LA���B�Z�! �1&�J�<��#D�	r���{E�)IT�q�\��^�D��ȠE��j^}�A*�1A����0pvar�n�Q�4��˜��_��M���� j���ƨX�!�Di
n'��smH�U�d��-�!���}f���_���9���	�1���D�q�� �1����_�;� ��u��.��y�W\m�9Y�"�K��ȃм�t��X��#�ʗ{Z���T���b���9���g鼋����q�%�"緥�i��{��!(����E���O/&k���I8�d"�����HMx��Ȱ�Z�iƢǽ�,�� 3�G�N��L�7M��^4�`�r��Mn%�A��y#�>���a���ĵ#��YM�U[��}�Bx���Ȉv��K�5���#<¿�3��Z"oG1�d������qx~�g8ڃ[��F�c�o�ucJ=�2I� ��7[æ)m�XlxVHYEB    fa00     3f0LN)��^D�$(�@�k��!@�o(�d���������㛸2f�iQG��'�5��>*"�n���UE�kB]^}�O&?��7V���.�����"I(�qQ��y)��ABU�����}�G-Ug�|���\Q����|M�P�?�o&1H���>���c{�u��hX/�{�j��s���e��`���{�m��Е�f��Yn1����Bc��8��)t�#� �@����w,*v;ȁ�f�@�H�놦I�\j+�X�8p�3h����^�O��L�T Sߤ*h������B��y�'0�b�3���x�}jy��]ƅ䈪��mx�>]Sa{}�z�KD�BI!)#�����������9~�wj�H�N��nx�M�u�~	�a��.^k��4�37���9����ޠU�.�r�<�T���m������S�����/������[;QN>��(�(�)�kI�����ț�Zp�%���Ѻe;q��4�V�`/m���|��͹Cz�H�%���ψ��=��Ԍ�'��w 釣B�=H�G�����K���n���?�����+8�F
h��Z$Exls�#���҆��u��t��~��r?�D�Z��\���!)T�E&�z�.�K���r5$���hI&1>����)�o���q�q��*tW�^#����T�E9�����eV��^Kl!���.�c�P0�lt��ܿp����h�M� �� ���n�a�P�]�=��J�����8ƕ� v{ۍ!H�2��$���I��h���G�P.Wtd#{�u����!f���DeB��)/��M��f�D�?����[��o�z��D������G��j�?��ߡ*�����A��0{0�������N�B��6ϭYO�\�ݐ������A�Ə��n:OO>�w�r� $L��<;���>��Ei��9_"��?A�;����»}����~b�d�}%u2�5���P4���Wj;��XlxVHYEB    8096     b20 MC���?%�]r�~$n����\z�Y�B&Nr��\�]���]5�Me�����^D�sw�V}�8 8tT�����F�v�5��PO���YR ��ٙ4�|�7���'�I}"{���1�e�l��Lm��� 7$��DJ��K)F�k%���8���=!Я�Hz���;U�8�M�GHv!+t�}�XQ#����*>��^��'hc��]=��J��X�K� ��}f����\��x�)��J��LP��������y+�R�׸�`$���
�GL�
j��+�W��pV8�1���gǊ_���gxՙ'vy���E%��K��d*���B8H��~���K���jy�c����H�0��Cc�I�_��O�~�&�D:8��R�Y��FoH�y�@L��|�<�"iKJB��-D�?���6�T\��*�C����ER��\z���R
%�Y0�	J<W���{l:��S H�9wZ�P,͔���\��.`�"nf4Ԗn~��Č��6ĵQ�"�ʃ|��R���Y�B</YR��À(%[ԇ����#� ��#�Q��������T���K�5��SXK]y�o m�DU�/g�ud�r�uJ�mj�qq��V1
�$X4�N�N�6����K����zU�#A�a��N�J��,�n|���DD+��.C+n��]���˱؈[�u��2�<�J�=���J���n�(M�fFXu ��T��&���D�.���"�W�$��C�"��i��'bP�O7bݑ���v���W����A�`A{����� �xY�ߡ�ln��y���2�]��Y랮� ]w�KB�-���%����e�Z���	Av�\���K�	�+�s	~��է��.�`��d�sGfDﾌ�~!����`��N���K1�����y��A�r��>!?ѭ��֣IX��L�D��0]5�V�&b�����
�h�3|�q��P�ԭ��E���0(D�%����dz�7���I�t��*[_�
[�-���V��;� N5i�98�w���LpD�e^������p��8J�p�L����/cT�WG����
�ZD�浂V�%��9����(�@���>}�/c;���~�'0���@�����rяԳ��B��MF׽Y��,͖>��y_Y;�����ՙ_%����7��������'����\E{�n H��C/ܲ`K��2�p>什Ja���7�b,ݞdr9����S�mj��6;����r�[d�ퟝ!��.�A,�?Dц��f9Sqob]Ew��p��_%��`�e�70Ҿ����9I�f4q�6���w�YL��#�;�G8�j�(��P�,w��ڡ],S�I�ջ1� E�Z}��^j��M��z��?*a�h�-)�yaN�������h���0���gx��&+���Qg0��>{���{u�K�ǠL��YUy&���`=�g�/I�u���:!M�UF��o˟��hf�����	���g�z/��K튁�x*��N��;���,��n�������J��@��;��OA�ii}R�y,�����_	�K��h|�^3�AF�!ACs��i��c[��i�-�ƣ�0�-���\������|�)��|��/�����F\�.;�o�^duGi~\f1���dզt�l�Ώ(�j�W�6��9%d�h���#X��v\b��bp�P�-��hC��6M��c�ɤm%�jQ����zL��z ���x"jn��!�Z�E��BS���〺s��/�� 8�����˻(<�J8���J��td����Ûo���`ʊ�p<CD��*W� ���FA�d���I���b��cnhD�8D��������쨹�l�W<��r�����*ާ�����+v"��x��#h���_��lO��5 �	5v�Q�)��nU�ƪU\��}�d�\1������G_�t����Þ/h8{��_�B�3�d��PØߏ}��S��=��#ϡW�r�ï�f�k�l�:���R#f�'��41�,���E���ߑ-y�7M��.lR(@r���#��ê��=�Mk#�j���y�fQ����6�s��;h�s���O�Oۺ��UT8{\���@]���n��YKx�O� ��q6
➳�W-�1
)hԯ[�g��R>�P�aZ����+�ޥ�Q��I?�R���b]*���6c��&�D�O
(��0aq�4�k=���υ@��s�P�ℾQ�lh��)0	�u�
8� {���հ�������eOm�:d �0���^���諦i��_w2FM��[�*J���{�]��<x���F�L��Eև��2���1���4�e��gaX%��G�*�9�&�1��E���Y�T[� �G�y�5��t�e�f?}M~�v�4݂C
�@U��6��#/t8�X`���D_�Zh�r��Q�`��ے�-G�������
9��A<�Lm.F��*�u��Y�C�#v��ni�)���u)�F��t����հp��z��{�-�ª��V(��pN�ɧ�-��Hx�Ϯ,�1�@�f_~h��1�P���Pfw V�XRm
��*W3$�N�X�239��z�u�t�e���8ZF�q�.-�w���J!��M�~�B��%!��E�,/H�<�pK�k�.u��Q���,����FI$��J�U~�6�����綔���E�5�z.\;w�Q.��G�KgO�h��$ރ�D(�L����7�e��2����E<�wB��W��D0��L:��	�l�&���:k��,?���@T�ImPS�}��5 ��Z}�J�M��w߭u_