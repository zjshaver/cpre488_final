XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��a�Ft���E���[qw���BH"���3s�i9RX9�>x�b�bmV�++C��u����,�%էc�!�ʷ��XE���c����B������e�(t��G�qKau��+�̃�%%��&��Gߴ��~GCX?-Ha���boX+2����ML
"�0���4r�%O�V<(F�^H�Q�J����m�H'Ȩ��gb�����H�}ܟ©��:�?;�����6�:������L�P|P��	Z����U��R�1/��fVީ���K�CF�XD�=�8��5�=��M#!�W���o���K���t3��sɅ��p�J��6��$����O˷F���Z�|e�H~1�pi�XH�m�������1�b�"N���A� ��8�ˋU�݀��ή���}f�ͱ�@&��Kg؝���
�#����T��]����-i&��E�h��OyK��1�h]X���m �pK���.h��,	/',�ˇ��-����>��ʓ߹��[�"��s�z~܌��<�kꦙ���|W=�8nuƷ��$�,�R)���N����q�~3d�_Q��������]���k0���$�=��-��u�o��N�@���< ��d�F�C��U�`%OAAt�n�$~���i�R@�Z��:(���I��sסئ��|v7+T-M���Z�e�P
�t�� RX�H��2���'���Ƣh_�{d߈��q�P�n	�@$����uǮ�W�"�)�i�r������� XlxVHYEB    893b    1e30��7&wX��W���"���Cہ�ō¬�hą&^/�ba�eXk�{|<�+�g�I�
[JD��u�0�y`���v����U�Kī��5�y�Տ�n�aJ���M��>�mӫ�#�����P�m�q��y����夕�wg�#��;�D�@xCg��R�7P7TMGl⬦y*zb��K���6������� n�D\|V��5 eu�����S�M5>>M�Yy�@�z*� L>��G��D����oׯ�4m���z	�"M�H�==���vO�Z{�e�#�
tV")�"����X~��ZZQ�ia8)����6��׺�%�5�����vㄈ��12� �'�­��%��W�}z�X�?hW��JF�b	��{͚��\$��+���ɐ�W'��@T����2��F�ܠme���|A��������Ņ�zԃ���hVz����{��d5�L�e�9-/\�dE��p�����;�4味[u+x9_D)'��s�1q�,� ���f������������T��p����A����%�hԍȇ�l\.	2�������	�*Q����B˙��{�Q�>֡gK�F�@6cc8b�xgŢ�:�iNo;�0@)����e��%e.X�W��z?�ꡏ_�ꪁ���]	�0��D���̖T��dgsH�#���foV���K����jD]�׬@�k#5����[�ܾ�X��5�F�ܸ��!aK�KJn�&V�\���~I�R��ov�3��w�gGӳA��w�pxaw�"7�9Fy�3�VVaB�k`�}#�Q�~EW���"���En��T�G����\�-����D�}��삀���I�d�!m(���OO?��D�s�Ҿ�^�8��Ƥ�E`6l����AݓE��J~Ut�9TMh`�M�S�.p�m��U>^�_����py8(����;%(=��r���������7l�Ұ:4Uwp���I�Ui;6$��FpT��Ii�1�6<[2���������DZ&៙s�Ja�NWC/��֬ټߩ_L~{��5���f̆%b�]@1���)�Yl~��|P��B�PS��U�%�L�S���;�9����֋��ܲ\��{����.k&������; d�T,��v�=��UX�	kA�Bhz؝�UtYg�5Nn�O��k](�Mז�����BA��V�Qw��r7c�oȱ��=��:�V����d�f��J=nM�VB�`1*!.�]�0�!?�T]�Ή�~�n�o'JNa` M�TN�Pl�[$��dM�'�هD�$�1tcl~S��-2^i�;�ţu\]�.Ys)�?+�Ļڇ�٥�Δ΅q$�s_0�Z��G�1�H$�Rd�e-��T=2����0��jԒ*�-��k�1�>�K#ז���M\�V����#$U�5�5�����-���h�s����7�� r�8P䟧��0{�1J�:�W*`��0)(�W0�E���o�)=��v6V�#��aǱ~z�� &Eed��$,b	���UR
j��$ C���_�~�;�pCO��/��L}�y������@��n���P(��(:���I��4Ɣ�MW�$�e��:?���c\�M���.��K��ŷ����W�l�����1�Ĺ�g��"#j�Ni�@K ���?L_uZ@�[ >*	Җv��?JM�j=^���`�~o�Έ���ػo�2�Cs3xqc�%�y|�f�\p�#�P��;Q/L��r�V"&��F����F:o6ِ��g�{���^�,�7�f>�8^n͌	A=����Y�\����l�a�"�f62��B���	�_�F����ˀgϗ��SdTt��j.Pi����S۟��|R�i�r���#mvξ�`�o���Ï�=oB��u�h�'۽(�<�
X�?�0��9_HoJMC���b����;ɘ�.l_s:Q�ڿrA���دED�d�'�;���/� �[ӡ�rC|_�=��R�'�_�B
����ԭ�Z/{� �z����4kj�����"%�A�N����ɮ���e��P��p�wV�Ĥ��W��L�?����4�ǔ7ᦫ� q	f�2
���#��:�AZ�x/j�J��%�[�3�$s]l~Z��P����89���v���V���z�0�+����D����+�0��Jɽ"?�G�jxb�z�?!��y;�2Ր��V�mN��g�$ʟ�����e5����b0m.P�TgN2x��N^��u�� t�cc�?����N��Ǡ#�2�J�[�y*���odki��!�NnpjF{I�xG�th����ض9�J=�eM�3��҈�|��q���\�j�;o��d��Z�#;��ݫ�-7�J��� ��uUZj�ے���w�x嗙���}ݘ����@�����sOI�8TL*k�㞈╋�>X�n;�UR۶���=T�	 �5��mX�����2��cp�d|
cS��Ah
ݸb�3}��-�x��J�lB��s��P��Q5l�0v�7�;.'T���h�c곐6�/�x�^���bwg!xg��hQ,5��8O2����Y���l��!Zb|�b#Bh'�?��<��4oH&��(�s��벴g��W �ڎ�VA�&��@�	R�-5�EVn�������a6qz�$�H�u�3^�����z1A�a��6���P��^t�Pq�s��Xx޻m�0�����X"��� A���}J�L�J����i�;�R ��1U���(x��r�w-��)x}0����Ĳ�:r��^8���p-��i�2�����!W^q;���+@P����I��Y5O7��m�D���U�X�J��*��-��L/�!7�H�#����yu][a��\@��cAa�����q���#/��#|�䮫��$��ư��_��F�ir��>q��v�w��C�9C�~sg��3>��|3�����Q�Y��c�P��qд��7,�@�l��d���k���o��n�/��2#���8B)'�3p�R�q����
A�|��Ų��6+��Պ����ͼI�W`��f7��!5�?���h�ˮF�A\��˃A]��mb�E�!͸ȟ0m.y4����*e-�ޱ�+%P���X=h
,��MD�Fx��Vx�2�݆Q���06�i�ؚ8��C|�X�d�h[0 iYT�Z��"��d^�!E���Zt+��>+= ���v�7���錠RG�r��l����\=��+������ϋ� ��E��6�A�J���;�����#��qu��N�&�;�k��ûhwF �Xw�ê��L;�����dR3HCj��o��Y�j�?�#~��#L�`c��غrޝ��q6�[D��5HÝ\���x�^�_թ��ؕ�_`%(�R/����
yn��!����K�H��v"�4�2�c)�aM��X�xh���n,6�hC��@�%>��J`����J��0.':��t�
V�ض'���}L��d۸��4b�	Y'���y��j,�QS|��� 	��ng�4�6�Ha�2\�O;�� QC�����s�������~�@$��!`m�jr����і��ۼ_��h�d�IC5K��֧rQߤf/f2�<��W+���tǡi��K�Lh!o�g��REؚ��s��C�/-2	��:�GI"�hr~M�����y鈉�����X�'� kGS�0ǐG�i��c��;�H���/�B��Q�t�����;I�^����撍��ks��Yp��;�w�HSLT��d\��v��h��N��h�	�4���l'�)/�"�\ME0�:¤C�~ ky%NJ��z�s�)<	�H/m�I��Z"r�O���m_3�2�b�N��(�b�jO�xľ3C^��Y���-Bl�	N�_
�7Y܊�s��<o�,B���}�oue.������#�^~	��\�(�֓f�U�P-�E��W,��FND��"Q�߅䀦0J�;7�;k[@�Mv2V�bb'�o�)c��� ���PP����y`U���.�D�b��B�}O;��(K3�0�|6By	Q3`�\�J��]^�7�$UP�l��w�{�b:�8w�M#�������Ђ�Ò��i���2��o��D�C�O��g�'��ݝSK�=�教͔<��Qw�a;��/+\ҙk'	d:-8;�d��$s/ԃ�����%�g�� ���|9�1�K�C4PJ$Yk�8f�c�n�Y��e*OTǔ�O
�L�Wl�-ĕ�%�Y�w^�Z�U՟K0STm
��N#�r����ܢ�z����k�2.!�2���y\eIFN�Iq�0�9m�+�@s���-)���G2��`�&6�/^��1?���Dx��xf��Z~ ?�L}1e��gq%����#B�Q]?���"mpt	��ݶ���� #]_�fa�6'���׎T���"��a��!x�+
n��M�;x��hJ�Y^��\�������V�M�U�����/(e�Ǭ�=>�͑ ��ML����(����~�sk��cr�׵z.Փ����?Vȉ��o�g�(�}w�]�>�ۖI���n�^p&�d.�vܲ(
M���X��N��x����	��w7E������8��6���OjT	1��O3�S��L���[�
@�2���A�8ሧ��\�bk�'j_����o��L�wz&�k�x��_ŭ�3z/��m4��U�Q>�b`�tB^�Ǔc��L�@|�6~[c3c4-ŗyh ����R�5��'���ݼt��;��љ�|�\�ܒof�(��c����>y�Aw��D��Y �8~���H4��7�Tb�
P2�����0�~�sI �̟��4�rI e��L	x$ZRf�;E���w�� J"�1%�5���#��%\�Zx}�5�2�i�tJl�� .տ��������ٯ?��E�{.b�("�����'}�̚++F������ϗ}1^N�oמ�~H�_c[����O,���%z����rN,*Q���e}��k�,�D�E��Ј=Ź`�s~�y[������*���MQ�/A
�����Y��k���S�B�� �8p."�zJM*koE�w�fŞ��|Lr.���E��~�h�#T	:�8�i[������v��=�D��<lϕ	cLt�
�b�cNi�Dzk���>��7ߦ_n�!�^����n0Lq_}5�ݝ��v�9j=zR?�J�C��p�4�o�k�_�	�Ēv���:�:�I������2Y�l6\���8f��3S�wzV��s�g�s�e���B�����AC���|ˊ"]�^U$�u��@��ߘ5��RT�/�r��%�9_A�0�^K�D:_�0c%+Y��+M��3�_�Ƕ_���[�x�=��e�zޏ����T�������gUntq���X��ɔ����#EOjs���JQ��.;�X+�%�;	��f���R{���[�9��D�7�7F���ؙ�&�	lF���s�v�������-0�[\��������?��a9gTK'r�E�'|^�|���{��{�ȠC�v��-(���yF�S�;�x����ӝ�D�۳�Yj��d38�3��8ڭ�ؓnE�d��5	�7�۲/�,��=�G�<Ζ�0�ձ�;�����Dl��ys����Y�G12�pP���M�^>;��6J��o�*|�P����t�E]Y~�'�V�{y��p:��G\-:B

=��	7�=�p�Vץ�{"'O�q��?=Sz�=�i���%��|L:l��窡ip���<�j[�3 �s��{�.z"EXd9�h��V�~�I��jU��T�ښ��d莵�r�y5�:������V�$�"�q�l<u���f[���2� f*
�pT�� �s���8��m��BgNC�GH�x�f����Ɛn1�S:-����K�|J�J�̅�O'}�����/#���VYx��'b#�'?e�@h�-#m���%�A�_Ͷ�.{E����}b������Ō*�����**���\uz��0f�W0�EN�ܨ?�5��R�#1����J�x��a�x�����I����\���D�����X�ij��Ϻj&��A.π�QZ_$\�DTڡrF�N3�����bN{�yGdq�Q=Ή y�a%�Kk�UƳpwU�L�:�7�(_N�_��������Ȅu�'�������7��\H�y�Qm/�G�����2�����l��W�����@�ZU_v�I{�0���}��v�90]��Q�E��A��ٱ���[��@[���(���Mj1�����%Ek�l���wݢ_4S�5=c&54d���HL]�[\nq�i)"|��k��xdY�o[��2Mq��%*�7�s&o������ 6�4z7g����$�-����uT�Q%z�Q�Q�uᶐ��Hv^�'jՓ:�o1	�W��qН��i��BX�_�Bˡ�i"��M �I1�z>��=fi�m��s-������֓/��W���1��{��Hn����ü��״���4�t�����l!J�!b��y�(]�3�m��)�[�����ܞ~�\l!da�'�u$V9�{*��l��7"y�[��6껜�覼�ZOTr���ю٬�vtzu��1[2�u�Ȋ����e-�_�^�к�	%5�p�)j0T�[gC��*����4FO��ċ5C�`�Ҝ�ə�ᓵ�<�S�֪�f�y�G��u�[*�8:s�� B{�䣴�c�aB8�rn��ɷ����9�o�C�0}���OdL��ߦ-V�38��V�SOr�U�W:�(>U���4�����޳�i�D	 ͍���&�r)�VT�Gωw�A�	D�
U�9���۰C�j0�ǿ���}Bf�C��XXM�B>�&Sy֟��׸ʲ�{�S�\U��s䅛�c6�]��b��Z3ͽ)�l n"M��	0�q觴*g˙�_K�]��б�Z�t3�`.�,������8OFU"p�����f5�k�fC`{�
��Y��l���c�tjV�O&:gSD�*\���-�G�.C.Q̤%
��/���ʃ�<�����T�X=�{���?~�ic��:�, �̎I�y�,�����pZ�7�@Q�k5����Ѫ8�����Z���̅^C<1�҉ ���	�L���ĝKU'��"�r	�S}��U����4n���Y"E�v��Q��+Q�Td���b[^~��⩉�MIV����3�e���5.2NP��X�:D�s�=�(�$l�ҳ0�"1^L��� �[��p;��ǩ�[ R��qbv#�ˍ~5%j![#bG�a埂�?���
^ƽ�W�ȉy
.R��V�C�2�^����_!@����p��mm���*��$��m��Ŭ�e�a���L;٢ę{���m�c�O�b��9����/5�;?B�_c�C��k��A���͹2h�!�37�C1�C���m�������"&��XTc#����f�[�L�E��Mo�G9�h0u�xc|Or��B�qEl��q4�w�2��?��x����IpT�Ld��pz�1��3[9K��N�	�e��Z�vtv��y��5�� �����M�z�������78E9:���j��3���nIQ<��f�J	B��{�l9�B���"9�LA�_�7��{���+Y.��b"��1���I8{)Da,.W����T�eර����=B!Y��C�ߨ