XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���}q���nS/���$h��Ψ�}>7�{�_�>L2�1��/�ohU+�|@��n�0uMBx��Rî�a������e{��ᜒ=�.�#>U�o�n=V����������!
��K�6�h������x�w>�M�M��&�צ��ɢ
����]*!�+X�_��+�O�N���/�-=pǝ�_�~�!6)���.��8x���t��I�Tz��_#�b�x�,&�y��7��W]�ָCOR��0��"��#�$�W��`����/��ʠ�}��1�u����`?=��7?�e}D#X��*h7yx�,��R�y�����E
���0ݕ)���N�e���[J\PP{2��?W.�tH��2�<�w�U���Q��� �#:i�N��7&Q�:;�b�ݧ�d��1�s�?ۓ�G�2�t�R����H��qب�P��>���%��z 0۟�$D�!ae�I�Ec��%x�"���~�nq�s����-�5�ؚ�������4(�4�k����P���H@<;]��0c�&���Bw�W2�!a7<T��B����*���'F<L x�=I����})[�Ў���Z����Đ�9mM�­t��	Q�?�d�_�:0(������ٲ���G$3�ͱ���'{��Jb^K���_㯋'�r1	���^�m]���MJ�^�¾����1|���9�ne{���(\�m��X�n��PC�%��{���5�m�Rp�vq|����ol?+��ڎ&XjLPS
�B&Jf�Z�Щ�V�VK��P��o��XlxVHYEB    1e3a     a20 #��ĦЁ�oc��h�_z��]��$b�?>K�<�HQw4$�o1���C�}�<�s
��J�.Co���5�_�k~o����[ִ<G����K� �,0Y�.2�t}�.�����?DD�$�SB�#�E�r�%���ƿ`������&�k�j�`��w&֤,����}	�y�ru�E�z�4����p	�#zZNTQe���ehKJ�Zԏ�x�Ya���Y�'b����O�l�JS�2?m?����&���4�D����#�>���ɰ7}|oB�D��>���s���>�p�M�V�a߉�A�D���4��b���|b�Պ�W���Am�*����I!�sKS+Z�a^<B�}=N����z&�{�v^k�?��I�� ȏ��_0�%�h!��@��0��V_�ӆ��G�B���a`8�ꉤ7�ى]��1<y���A耸r���tf�%�/�{��rX!����m���!3���vn�Ж��]���.�f[�0����C�Y���2�c����a���� Ol۝՘MB4ϰW��n���
.uuE�Q6`�]��zJAygߚ�m^͢~����CU6ݫ:��:]z�I@Sh�W���9���V.ń?H�9\v_����n�~���Cn����`z;�R8dg��l_l�O�������0��:��7����)J��пФFRY87E��ّ�VLD*�V�5w�R��"wl��rH��}�;���L�ƪζ�P1�b�Y�{�,��r����,������j��{I���P]���Ф4Ǉ��i��G��۳Q;����S�5N�-������'�C{�-X����{�s ��^�4�'�2@�ޠ��7/��v�Pe!���
F��9o�.�X{'n��f�XagZ���+2R�3���^<D�1�
	YK"3���V�E�TB��_3��Kv3_�%�ұ�� ;��}���AT��R�~l����Ĵ�fh�U�>��&$�����3Sݏ�'|g�>en*�o�ơ;E}�F^`�'�o�������.x��ʤ�g���R^{���	=`�1Vf�%>�,	�	�)���^���5�G`b5���4)xՅ�αy���!�4��(˔�1P�h�͜a��������S6�U��7�H�	����$K�
�r)O�⤆��2_��Im�4��z*c+����O���9��^we�B�!���R���_������{T�'�P��w���*�0#�c���3�1���E(i[��| �hڿ�7���zN���xxg#"�GUA)g�M>S>�9x=`e6����1�ٔC����s��)p�s6�DU�**5�k�A#���HG��1z��(��Q�zO�'�q�E)�<�%0��f�U�CW�v�Ź��K])���P!1�j�G��"LX�~7���r4��:|�ӭdpRg88���Ft�?պ�$,�:H5BxjŻ�cG�AB���~9	W��%�>!��>N��S�ek�I��~�a?}���>ȹf
{u8�~���r⏺Z��f��L?�����E���@�s��+t�{8Ը �CJ�tiA�.oۜ3�g�4R[�?%m�~@�S#��͡�і���Gㄈy�]���!D�z�J��}F����F�l���5�y�?v�Z�J��BE�2�B�~�2��"?h"�u��v�����p�~/��o�؋�-�O�J�.Y#mӟ�U3���yx�D�����V�脩]ˮ?��5�@[��T�)�a��k�^I����~*k=�9�f�ShjUJ*�e\U!r���@ru�r�J��S̾�s�I: i��-GV� m��$�
��f���}`Od�b��<����41�]��Nu���D��4Yz�H!Z�g�ښ´f�T*u�����X�ځ�I����f�4��Kg���A���n��i{�7��͐�e�#�?F�;t�:����D̡>ZV�#�s������Az�]�|�W���&uB��)a���E�¬_"��1���G@Y�U�Z����	`aYMu$�L���d'��6�{���cѸ���L���/E����|G����>Y�T��q�n��5֎���Q�B��&	�U�g%{��y�����S�%�d[;#CV!>�`GE��RA�o���.٢��0�[��p�� �����M"]q������g2�v׸{��1i�����O��U���,��{TI
��u#R�Eo|��K�՛�e����&��n�	���� ���5̪g�j��c�瘌�K��T���:�?z_���l�n�z�)ڻ�j%��
)�T=�p��{�\�n���62��ޠQ͹P�dv`�F��N?�5�!�+�$���T�\��[���i�E��H��Y���Y�ޛW.���'�V����:�Pv~����L��"�N⬿�/ګ��q�_dC���6�W�S۝�3c֢���nw�� V��z0ȩƖ�Ya����L��X
�L�1j����-ݿ�����!��mOźsȵF������?ݪ�; Ǖ���qr�X[�4�7�ȏ[�����ر����+�-�V��N`
���,_��iH���Y3�