XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��1H/B.�킧"����b�ŏ��J�<2+e �SK�1�]�"`��l7��=q2B��
%�C��h>d��2�<���'��6�1t���wt�H:d[����>L��T9����}���ӆ��	��N<�ʉ��Ag�6.�]�������$�l��Km,:��T#�� ez<Ǎ�� ��"�!%���Z��;����cP�Y`w��G���"U�s*��Pj��S�;&��&Nb̟S͊0�Ģ���+�{���N��N�V �;ZC���|��y��sG�S���aE��sn���<^��1p\��R)�y��� �ʩְ����e���.D��?ߟ�.�%��m8��5)K�i~���ӎ��{�� �1W<�c���g���7��t��n�*X*u\��{aެҮ�cJ���!�'XWA���hw�m8{��@Zxgh��XdT�Y�C�4���9 �9 �i�~XOzV���J��G��
x���7?���C��؏�[y�v00C������bw-:��P˱�2�H���{��8QF�=h��b8��e)h�)������(B5�VA��a�>r;�_��w��[��]Z�V��V�9���MN����<F�6������-5�_%�*�ii��_�`m��m�s�.��,�����<����W O��2���n�܊R�äI�%�~E�#���=���l	|�3d.�t�OZ�7��V_b���zO1��T������V��	i���PT}ߟ��u��X��D�8�:XlxVHYEB    15b2     890X5A�+��Ҧ;[�LΞ3Ɇ���c��������qY��Z��)#E��RY]��cX}��V���R��*�}�9�^d�,��piMMPs-���۸c���KJ����7iaԹ���w�é�z	�}���`*�Zւ����.OP����jo^�V�lD=ʥ�aAtҡ9�`��!`N�__���O�I�AA�Z#?h��<���C�G/)ϯ�2#���<p��;=�t</G�����nD���.k�� 6be��_���?��;����ͷ�j�|nɨ����V�̖GZ���DkpS[(����9c�����x�r �i��oY�%	���OC�ʘ�g��K���(0He�b7�W%k�R���'�� L��=�I6`�(Y�k�|fb���U�Ip�"K���#) 1���q�+GiE�b/�����k�� ~v��h�7�"[R��do�;�A:���>3����:z��mq�N����e���
�_&�X	"Ӛ�U5K�^~����1���97�LųB�Fl7�6�0�|V�3ݧ�XÄ�r8����{�1� �pp�G���ƶ�V���IH�1U��xTm��z�	�yKx��9�����l���V����vk{���"	[,i�op݉�������+
#[��;�M��c�)�$���,"	��]�h5�U�b��6ǜ��_�/���R��R/�Dg�渄��x��ؕ�!����� N#�ef�X4��E�
�k��k����U%#K�wՐm�=�$���/�D���f�ך��/T��i�[CĘ���a�e��x�4¬swL�LCc%g�r�����	"�5ц��������Ƭ�����2�SM]�u4�V�����;���$O�$I��pS��F�5��αU/=6�1�ǈ�m�l����1n��_H�IQ�#f�D-e���"��5�t��҈C���mZeYRlOz�s�Dib�o��#4��	z�%Ï�~ O8��	�br����{��HfLZ�GuhL�3�&�
�����y6����2����R������Գ�&��Te\&VX�H���k�ֺ�'��A���h�3
��3�:��ؾ\߉w�h�~��4�[���4yX�T����wn���y�mx�/X1c��Q�ۺWv�N�br#��x�����M���f��y�r�tAcYTH�_u�)]N��FH��2RE&��7f�}�I{pJ>�RrG~w��R0��;h��?=�
 Y+'uWnM���[�ғ��GN@����{B68���f�b��M�kݩ�0:8�$!�~���'��+w�뿤�(!#��������a�u����(a,�)(�Hy��L�}WP2d�����n�&�/�>'?����qX���Ck�y���것7����U�kl�vr�Y�����?��j�oY�
E��[ӴK���<����b�|B��b>�O���{'���Gk{򹥁�p�=��j��k����B�pv�� y4jH�#M3�ٽa�T�0���C9n܅�6>�Ȱ�����\�ߔ���6�ܯp(4�!�\�����j
����
�����!ܾ�(ί��h�J�T�o᧦�Uh ����%
p�U�,s-oB��ݥB���@4��E^������^��z�Q��&_�xi(R2U������^�-�|��,#��š�28�)��MV����#H �ʺ��敮����h#�����������(Bt�<��u��k�va/S/���2�#�.�C�ŹSY�g/��|�I� ܂R5�r��[��|4�N�(x˝�ND+��)��́�+�D�M/�f���׏�H�=�����$^�M�b0�}ov�`D�_g��J�ԶM^d�g�LԾCot�axֲO�̑�Ȫ�bQ��[2K�A���rQ/��H�QR;`?��L�#��x۳Xƚ��Kz<�>��ǫ��p5��;�ΰ�
����%�F^��F�0���N�#���{I�ҕ�	��J��f����"Æ;[,��D����;Qd>�=fʴ�7>�g�	�j �]ʏ�3�"��U��?�O�!7Oh]������E���bK�Jc$��q� ���lP��Dnw�+�v�T�Vf�2��)zY��R��Ε�ЉkFT�k��������j�"�I�U