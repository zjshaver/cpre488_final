XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��s��G�A\�k���^K�L����W���2D�Y�T|M��KD��ذ�Zu�%?O�,V��K1�^��0⍒ͶE�5P��R����W}+��7-��
�(��3�ǥ-��"�!d|�I��,�v�%ݐ� PTc�f�h�3�tZCU���5�	{��Mx��")�-Q����\9�iBb�����CZ��#T�'�ah���c�P�Iu�(L�V:r�y)ZN��W�3K8��I0ph�m���F�#%�k;����d����Z�K�M�i+�_d,O���.��Y��#�fe�no��?�%�@����ʜ&�BN���w<l��~�*���O�@ao�i�1��?|��Z,ť*��讆��h_f��8�=x���:��=�j�W$���/o|8J����y�_ _�X�lzZ���E�.����.�}5ϔ�6������(`�M���������-�n�MpP'Wȴ�@�n�
�ƾ�R�iI�sZ�--�d�#���Y��71\l�>}��0��(���M l�U�I�������ϵ�/����^��C�U�7�t0E�ZiE	�D���4m~t��煉�`�_�o.	\!�xW���ݺ�H��m����݁��q��k���Y�G�)J6�;=M��H�f����bԉE��Ǯ�:�J��%�{�;�5�Y��h��N'��ţ���N�O�OlO!Oi#���n��E4�f�NF�[�(�my
9)/ol�H{�z�~�.uOR�&}�����\N�(B�XlxVHYEB    3fdc    1160;P3B���5�_*p�O�IYk�ܠ˱��[��(RT���4_�s�5���T�
��IzZ�uT�N"��&�<u0'fi�y�6�$Pu8h��s�'���$�5��u&&{(�ge2��{�.����b�KB�O���e�>9{�,�ePSfǂh{�Cud&K�����W�Ib@5���#7{t1����y�9o�V�ț���1��_��N�7����ߥ#\���Jɠ��=��kÂb�q�k�����U�Ǽ�l�=�A�,9�����C*e�6��VGM���hq,V��ׅ��z�ꤘɯtQ�B�&��$09Ai&+(F�*��?�¦5������xȹ��>���x٭u�L��5H!/�,G�M]9��5�����9��\>&{�Z�&���F?>1���&E5��p�A?�����Ӈ�Oq��Gj�kX�ݪ@?�8�P��1��-���d�Nfv\�Z^��E������J�pY��h�b��!Vj�l�;�M�oh�S'��� ��bG�0JLl��[�;�nW�% g��,A�8���鋶�ا�@�<i\���N�H�*���nn7����7��}R�V;�Q�=�Bh'I�b��{����=(�Tf(�eicƛ�WM3���@g�1hg�7�qI��*Q�j'����S�y��N�6=���OQs��8>@~�s]VY�O��	a^zc�.UԆ���U�f+������VR��q)ehfe�6E��?�R�S�����*m`��/�������bpTJ�����]�?A�$t;��Ϊ!!j�چ >f�ؼZ0�N��*4�έ�+�s<�ODn���+9�:z���c�T��Y�P($�5�A�Ʈ�g�K9J��<�a#��"�O^��sr�mr�2�n�y'��˪�r.�u@���F	/Pܨ7��$�b�
x�I��؈>�Nl��? i
wL��Л�kܩ����Zs�a�F�{��@����39��j��q�h���P��S`�<ʙ�{�b�^�CXG9)ӳ'�L��蘌磙knIi.���P��C�A�k��5����b����4wU�e��� �ǣ�@�Q�@����<w��7`b�݈-����见���%�ݘ�q�0�ۄl��bܲ�8
5'O(KV�G��g�zr��ꌙ5p�撵�4���'��S��,]�0�p���qQ����U颐�lj��<����n��l2��,�\a���*����FD���i_��o+��3V��Vk�r����)h̦��G
��	{�|Ͷ/?ւ�caY��G�
�-�L�kR粚h�����1*�X
�3⹖�`|��S�ݗ�=em+&q�f�X;�M��<0�+�y��]�hq��A�
�m�^����/5,[�o��,v-[��c�#d�Hr�F��?4�����uj�rk�9�4�?L���h_���� �TP!�-�D���s��ߠ޳�^�&���<ncn"bnfz�G��f�@��)˿aZH�߿���\˖9���ܾ�w�1�)S1����AӟA憭ҸfC
P����䈍?[��˚s�H-�ދ��{w7���}�v,%\��RU���t�bx�%T)hVز.�f�ᩓ�g-WxO�_��6l��@3]�b�[�߂Œ���PH][A��t�<.�x1��g�/��H-�g�����qV <���i_��m�[���{�Q)'�
D��!+�����$���F�=�i�r�ʆЗK�?��E�p��6<"��E�88$�?t}j�:���|���e?���_���ŹCF�U�-�ME5���z��4L�m��Zܡ]L\8�7Ӂ�>�Y޳�.Ȕ���D��f��2�F,�H��L���^7@�M��i72���y<?�Z�?�-9(��WqPC��ϟ�a�'X߮6��f%+�]l��ɹ]�4l��_�bWR���b�~>?��-^�>l��!��VB��B�o���XsUrcv�9��������!W�L.�?q��Բ��,Y�L9�	�7L�;G�`E��5Wڎ��I$S#m�����ӄ���C�餥A��P��[m3lL����o�ѴbZi#|\�c���{�	��3�ʫGR�qf*����Bp�,�r�)Uሕ�cjD����p{�Fel���X�]������օ�0�H�%�i�]\%���.���,�Y=T9����u�Ԡ��Q۰��}�lU8Z�@T�Wi�m	D�X�f9�� J�,�+�c
�� ge�x�
>�1�f���:�o�u��4ȇ}�5����_�*�[��"v�'%K�J���C�Y�,1�|<y�>���(��ǒr�4=��۠B�J�f띟K��R�$���^��0`��"Lf��8�;�G$�c⟝d�����r<�2�*O��,'[c�x����Fɖ[���<  �����BD�M��'�_�z7��h<�-�x�˵!4�� �.˝����l�*=1I�s�]i�{���w??.���c�v,z*y�8j���}��{�ݺ�Ǖ�g�h�� %b�v�,� ��PW��S�u)	�b��>S" �j�j]�d�z����z?V���w�P�I�[fC�V�y��dRVr��!�5s@Yb?����"Ӫ�V�g�f���`-~�o�� � kXDx���(�X�ӕv�1�L��suۿؿ8&������S�!�H���Q�c���B����J���<@��!����H�<~�so�|1���C] �޾���ⵜ��Ī8^���qƔ�4�ͳ�nn���7�g�D�;!���`�o������A�Vٞ6s��y�rqw'�m?������4�T0ZqL�6�8��;�Чҟ��#�y2�=����aF���8�<��2tͣ6<X͕�� ȓ"��������m�?�z�<c��w]�{{�"v�N�b�J�M"Djeu�5��	,�0.K���B�Sc�m;��l2��b��y/yb8�E2t��ǎ{��	���?;[����H���^�#�?8�c/l�VUj
W��6�A�9)�R;�v"��Մ(��Y٭KG�P.b8Ǫ>�׺�4% ��E���\Tc�]����������4)�F������L$?����3�,o��`��ڎ��G I{�տcw����uz��G��
-��tF�(/����:oim�v�	j�L�_��
5\ҧ�ޏ��n8��9�����V���X���$���8O�r�dY쐨q�hqR�|�m�ں�H�����9�Ci���+��������.��}�Ӎ�v1��Ɉt�#�U��ɇ��M=t�������jl��������Ŗ�)ꕵϫ�j�� Q´˵mt���W�.KC�n�:ŏ�pw��8�ꘚ��C�f�J�04ΥRfV������}�az��Z��#��1�+A�g�j�V���2,@(�b�F��I..>��U�&$r�l/ڑ%�����˦����L��x `2�����6��2�jӬ������}�Vd����~��0�x1ؖW���V�i8O_:Ym������y8\��*�5�N�\�h;�����ɳ�ȍ7$��O�(ڼ��C�6�-��L��Rf3ڲ�#L���K����J���!�+�����S�2�'��`%7,6�B�Uu;�yE+�% ��Ab��]?��Fd�+ү�䗋Į�����}���s ��Zl'� �T�f�r斊(	թ�$0�U�bh�R���?������b������)�?!�Xv(�fA��;�r��T�x�z�@GW��F�Y��˨�8��bW,�d�r���s��G�FG(E�ޜޔ�c!rro��N�ʸQ�t���#��u���"����Mz����q��e��nW�`M�J�$]�@� ��C�ۘ��"�������>��}L:��)S��c�r�Y�Z�u��#�uP1�F\ۗS�H[�d�m{�V���g��L�`}�aU��V�7UpH���m�Á�h�I̶W"���mIk��;25��AG�YT��OfO�'�exjgV�R�ϡ
>���(�	��}���&�i�S�h!��`H�VR$5�R`�I-��!=!�-g�'5M'u{��YǏ�ȏs���n��y\�y\=�V09(@y6_FY��o�>�+-�*,���[�f'�9��O���"�����lt���V�H���L��D��˵�G�da�R^4�<o}e��0�J��P)�v�:�΂������7N>5����N�Lm����	e�N����ֿ�AI���,L���Ko<��̀b��Ԋ��c萧�&�y�3��#�\ts���Ǒ���]o�p-탠�T5�J���^nY����,d9�&�3�T�� ۂ���Ԣ�U0ck���EǷ�n�z¨��𠑾t5}�&�i���ִyXP��B�����y,O�-�h