XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��f��yx�M���#�Qr�f,��&\�8� m����K��U~��~��i�h���*2<�S��LV��z<E����֛��S�U�K�GK9�>��}���:{���7�ӊD� R�JIB5��5��|f���f,�=��ަ�FR���V��y��n�����5J��� l�`V� ��k��GJ��{����Aa�*��$���i�h>|�P��'%��a���T̀�7��AM�<Xf��ད��452���	�r�%ưCd��"�[�IG�Y����k�'�3�έ�bs'xOa`�P���1�-�y��lR�_�Opm�c�g8
 U��f������?o;7/'V�vZ{���V��׫�����9�yqf�v�<�X��-�q&�"�C���{J`��$�K0QB*#��7�_�:�>a��H5��m���f(w'h)I�ю��|����G��
���B�������+}s`�Y}m������;w��(���-28?ڠ��KN8��F(�^TY}��f/T�|����܇;�Qd�B#���G����䁘m�E��Y�2!<�Pazq��CDR i�6*)�i��j�n7$;^6h�ȺJrF>�KR�TΞ���u�kI���B�s.)�3��/�>��^Mˬ�^\�:d����_ۍ[�V��}�p�Zzsi>�-�k�;o�>�'?ܫ�PړRv��RQ�q���N��S�0(wqm5��Ө��k}���e?Z�"-6�2<���2��'�>�u
M�XlxVHYEB    1ea4     920��?���&s�1�S�q	o�i���#|���E�r/*j�\z>�|\�v.Ҫ�'5�ް�NBd.�%�JV��e9 ׾Z��4&Š噛��.��Z�R{S{욎��������Pk��(z5)��P�����Lǹ�?�J�����n�/������G$���",Q����<�lO^�CX��TS1X!d _C�$	ǌ�M�▕�˿�}Ml�/�2fJ��x�oj|�B����3/�<�|���>�X�_amF�h��JlK�Xo��>���pk�KX|W-��v�p���'Qq��̶�[���E��ڊG�e��pH�U~lD���k3��;�/��[%ZHC�Qqg�OO{���5�PKw�A*|~OsuM�]���nzfz��ծf�t�~r7�~�C���A�b5����I�|�3�������ۖ!N�q
p� EV���|I8���
�+���c<��sHœ�?�ܔ���M/e �u�\�F6%��ަw�i�|�� �x{p�ͪ��[�Y]�9+�`BQH�[u|�n�+)t��X�vԑ�`�bo�<�}7���¦����d|��-�^���]��&z@"eG�.���v���>���E�
�4�	�QW��a��1׆æ����TqT�=�|�"_}�*��nh���-�t;��i}��8�Y�Z).��װ����`�`V`�k�7����W����\�mi��!��y�*�� �$`fx�zq�֩6�V�ib�O�ȟ6	��������6`��$m�Ȩ����A@���[B����8�Ei���C�����!$"?��Bf��7�{�Gb���vЭ�}��.d����h�K�-�Z���K�i����8��j��7��f��2}+�.�4ct�����޼p+m�ј�Y{O�"��廟��2�!�������[�4^�7��7�}��鮃'X5�}$����wHN+o�t��J
n��c��\��������g%�nU@���Dmb]FZk���D"�#,���<�f9�!�N����86�ʨ��k6�ٻ%��fȰ���`��W�?鸆{�yl Mǳ� )K�K���D
���9/j���^%.�r�4��p��d�#[�F�X����?�]�'�~�j��>o�h�h��Q;�]���pr`/(y�I�j_�[-����\���6�(�(��3Z�s�/ߏ�]�V�0��_���{�T<���O畃�b�g::�\#I�S������H0��/�����5UBf�v�'e���C��>���5�Ś��:;�l~�@F6���U���PH��0PZ��y�1�(',ͣ��t���/��)=m؏,���\S �V�\���s�u!�����b�=	�<�~�>g4B׋��O$�&�����  J����<�b����"���o2���O������Z�f��^s�;�	��:�e:�
!�f�7"󺖢�0��3>㻺8F�������'#of+�h��9�|����������<�ա��(l���ژ;�Xmȧ��K6{q���xg�����������)����^F�?Z��#$�)Ν���H�iג���1%�&m���d�.�����f�g�)��8d���*+��蟸&\����>˓����:ࡸ�6:D�*�,Z>~M��¦��6�ϕ2t#����<�w���s����)��~����á�(U�ى����B)3-1���^d��_�#49ςO��^����T(%@�D�Pɲ��ԝ���m�#��3Z؋�H�Nn�N\�A�E9������%`�D���>�IϨ^wsס[��7qbc	٪�i��<�F�ξ��Nh��9��;���!���M��N���,h�ż�W���/ Z���|��
�?G���b�m�,:m(�՘mA	_q)A9�!#Xqb��Bt�`��$_����� ��Q"��M�������]B�A�nT��<��aW��}D��Ƕ�)���.!��{�9����A�퇭w�}ځU��+%�4�;�^Y�Qђ��{e��'��1"Š��sY���{e��L/�`��������S�5�zdYе�A���lYs� ���k�x��]w��?���n�C��_����Q����Ӂ��Ǩs�}�Jg���
�XS0"�J��}0p��e7�᯸NL�_[5�勘ҧ�)f?v�e>.W��|K���6_�� �9j�-e�'�34O<��(j&ͺD�4d��	�k7��Js�&�☹hLñ�.4U��Ʃۢ����'��F;>�8��	Z�kV��	ďz(S;�L(a����