XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ya i�ͩ��K��r�]��*��k�g��ӡҐ������^�2sc1�Ɂ3��^_����'���X��}B��$Qh;�tl�O}����}ݺ��Ek!7�RP�+��4C�0�$����ͩ2v��:}}�&ɼ�H������2m�&aa�c>��"'������]�j�W#�����Ob�-4s~r�v��G^�&���j�y��j��:~A��(���BO���ް&��e��o��m���P�x��P��_lt�D�0@L\rY4)G�12��`<
�,�@���OH�F(��cTN���F�˦�(h#R�����?��ʖH`�{�0|�;�an���6[�F��wgnc�	���jD$��b��t\�QZ�d?f_s`+ؗ���a�+s"F�z]�k����i�2MU�d2��k�!E9�Hߦ�Ey�F��	3ukye�<z
2D�b���2 �Ll��S��<R��?#��	���&�w1�	�7F��.z����y�V4�V�*��k���\d侜��K0�n�|I�S��(��V��L�yn �i�n����g���퐄Jng�y���t���|�v�W�Zk���X�x�ǫ�����x���㉟���Jړ3]�y�k���~�>����Lŵ�U�⴮a���e�����p�H�ER��S��=�i���$~���'Q|tb0���ؚ����� �8��X-ƌ�ր
�TP �Ծ��W����{�s\��2�Z���[��Q��"{����>�?bE��Y�nB؄D�L����XlxVHYEB    17b2     880�5��-ǿ��߷M^q�
�Ue `)P\z�U���n���Ԛ�}@Y���u-��v��zi ��t`r0� F�����C� SoTVg��A0j#�s�i�i���JvfG�[}3�׮vJ{�FJZFw��Af��rR��K�6�_�
,_���}��Fw�1G�M_�G�6�+T�l�����~��k� �����c4q~hWڼ�&���ĀY͒4.o�����4��Q�ݟ�����U"4T��X9�Kr��i��� �+�����.NF��5�sK+�t����݄����_禴���3DX3�{����u���(��6m$w����#��88�F���~ɈJ�q��& �j�#^������o#-�ed�����!8W:���1h���4��v�YLSJ9E��W1i�.~"���@��@]b�FZ�K���G�&�*�G	:�ðv'����G��gP��� ��P�V9(����[�l���Y#u��FO*�!R�~ī����dƯ�t0�c�?�6�$n����X����` ��J�c��][ڡ�H;U�U��j��A��6A�x/J"���Iϗ_���G��<�q,��O?�_�R�Mǯ����u�A:�,#�q�G�p5����̟��Ͽ�m��-ހ�UO�m_7�.���=�zT�Y���!�����F�?N=���˼�#�J���KW�	��S�X�&�$��QQ���l�K�����~Q��(�e)Ď��u���+��қ�}7^���7T��gz��᩾c�?	Ҙ��UOɴI)��-�=x���~{!l=�a�AJ�o7�a�����V-����n`���S�������~��6�Ʈɬ�K�<�ᇎ{ź���|#J��4v�م��Ӭ㑮)Ox�Z{/gP���}"6h _A���ޗ���F!�{���ɱ��B-�3�E�Z@���;+D��')u�}U��W���"f~�ޔ���}f���j7"��_b��F��I]� �+�wޠ��2�GK���k�Yo�����{����}jc=�g����i�Y�'���p@�\��om��@8g0���Ѳ��}�|�i����9y�T#<lT.�m��U@����I�-�A�������kg���4L��	1n�ڲ�S�:}b�3ԯ�1�b$$��fMS�KH�@�j��PE5T�t�6ݽ�6��y,� {oA9�E:�����FA�(����ȡ�n��߼�S3�B��NT_@�tF� �ރ�G����(�H�ʹ�&��5����h�����<��]�ju�dX�l��˼���o�Iw ��<U��Ơe:�)pK�c��
�p�������ژ+�C*k5s��u���]O����q���i?Ⱥ�-m��\��k#�g������u�^:�h�øNu�6�B����e|�n�.���2���aHrT��ՅRjP�i���#N�e_�Z.x�ѣ�s��e�}]R
�Q���0�$�X�����ދ5���r��$�ݘ�x|YJ������	 � о)��W�ls�J��emP��x|��+����9�F�6÷iw/n��h@��f#?�ˁ|��P
AM�]���ղG���(��=6����*'E�+��ve���7�D��8��fJ���
�O� �R��a�.�F0��>l�jѰ��QǍ��;����Y�����>R�fVξ}��JgZ-ԛ܆�5��0f�ū�=ݱ�,I�W(Q��Og�b~��vP2SLwt��P����+��N��}�yϧ�����ǲ�P���5y�A
�f^`����:����Z�5NX<c���f.�73������z���:2�\�I��S�V(�7�*�,={Yt�S/X��Sxêט�0��9����b��N#�`m��-��@���y���I�@�t���S�`7�K���.g��s�T<FK��$(-4��;��,?�[���@*���gu\��b������>a8U�]6��i�����@14��	��nļ�U�'��5x�9T(������vN�b����)�b�}&��'l]�K�;1�cPz��a�O�١�$�e���1Y��Q9�0�y$H��%�k�������4��RGl�c��;kiL�5a��w<s�s��g��b��8#�