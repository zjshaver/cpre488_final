XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���~�;d	��qw�Kɓ
�CE	EIX�e�'a���{���߮9�f�-8f.�����ݍN�Qlv(JC���Վ?������RJ<xO"�_<r^D�5�p�H2�O��B��)"�9�����i�j����w�nm`%}�q�j�����i][��5����B�,�3!��R�0��z�z�����.�m�)���6-�B��K��ŻQ�(���Ti��p� Y
�H�vh�7����Z���g�)��ޟ
d݆^`_�HO"�P������Ws(\�Dv�ghO�n~�s ��)p��8;|�cS eO|�g�k �nr��<S2�ܕ���J/�^���'nb�:�o�<�h� �ާ1��w�@�4P��D��x�1�DV��!��&l��tn���J���s�X�&C�3�)ֶ���ۼBcFzgn��6q��T���9<RCU�Y�B�<>�j���|f�
� �!���(��&Un+ώ���	I�L��ڻb��T+Ĝai,k��v]BgA#|N�h©J��m��d��л���KoRp<>�j�\^x��<a�3W�7j���]myN�鿯+r8�|�Mo�ߴ\�F��Z����5Hd{N_��=����#�@
>�vp�;���d08�i͞��r���7�, 1��]�S�#�R*^c�t�'��mU�¢~U�p������Z��`����K����-���=�ܞ�'��<G��q�� ��2˿��=M�`E�\XlxVHYEB    1448     800�1��Q��� n�zH�7TIX�o10��4_T*����֦c����Ir��[Y5	���u8if�@6���������;Őf}�8�h@�J@���ph? �R�T�>r�ke�ј��ՖY��c@Y���B��1��*��/��[�Bz�e� ��9�����/�)*3	xm*�����W��4)I#}��T[�Ү���(����B���w;���Rc���O*��b���A�-��(U�,�� �7��ZY����Z��E竓cym�M��ʿ�p��՜��,����Z1��&e�2qԎ�t1��|�N ���B��$���͖I��j �wby��4��c���Q���!a�"��)�Q�O�(&-AN���H�tEke��&mV��ٌf�e�9�ڝ�J�@f\�]��Z�n]���3r��cA�(��[����Ihq�~�������w���'}Gh]��J5%/7�՘X$ �4V&��^��]b�߻�J;1��G�h�v*�����9O��IHo�n��x������X�6�@��ӥ-M�����r!Ł���RJ���a��R�X����Є�Y	(I�H����"�Y�&�1buEuoTݬI��"+�j"��Ơk�C+��z}�d��3��(Qi�{�4�P��w �<�6\�0DD�>��=�����zby�or̍i?�bo��l}G�r���D����5���ٖ���TVzi�d0ˡq3��XY�v�]3#�׋V�?P� 	9E3����ƈ�l_M�s;1�G#�]����G��{8Yݎ2��	�JXH�l�t�)/Z�Y\�.��RDE�K�=�0H�148e.��6C��K��|�l�.|�13�����EɎ�4+�$н�fr����L#�V�]��wa,�x'��:���¶4�kP��(��c3�W	�8j�̊�PFo�y@�N�gD�&CY�d[ô���5�@?H���x��sF,�Z��1����}�&��N;�DE�����!1��ڼic�%y�)Ș0T��]j��b�%Φ�������W��V#8�~�R�����	#�^�h�ERk�PbY-�!�R��Cp�p�*��G2���Bʣ}�i�5��<�])
6�+ۘ��ݷP;W1-�7��!�0P�Қ����s�����B|=�����1'�"�b���t�5f'�1��HJ�ٵ��~y��I�F����ǲ�;��މ��c]�}�_�x0�7����'A7^׽����K[[g-�v����[���S�r��1\���G[����N�ja�c�XG�i�#/��>��L~� ��xҺ4���@t�g�O��A�gQ�l�#87X4��JJ�0�?RC��vP��뽕�`���٣_wL"�a���/��8�ϗ?�F;+|̭d߰�d� J����x�,��<��EZE潩:N��|V����j��Ҕ���p�X��,V��x������`%EР�2��^���x۸%���T�&�|��`�r������G�ֽ��`>�������<y!�v{K��o��LNBy4eI EP�fQ�<���@\���1��]�o�G���@�|\��dW~"�եF�%+XC��熃w%`����f��}�� �Qb��6zF���w��H>�|���h���6`�r�]��c�=�g�22�����Ļ��+����NU[��us$���;����}�|���b/͙��y"L�r9�/�3hݛ�9^$Ɂ{�^��,�>A$1��@���-.!��01: a� �=�4ʑ�X�|�˲�� o"e�@�9�+r�ev��BW�Q롍�F�U�9Շ8��T\:d���wP���>�%Q]+�.+��,�zQ��ȷ����� m]�|X�Z�?��܅��^{pX֏-0s���2�)]���LWE���'�9�M2k���k�������9��ڨr>�C䔒ؿ���8d�̯��5��:�	�.Bx4fHp`�C�f{��s���!� ߣo�XӋ����$u�����O�Ww�����kL���	�����*=�Mwe�TvV