XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��f)�6�攽K�o���毾$s�ѴH2����vhL�W5�1+�<؜w֟��Mu���R�l̖����]28Gc�t:�G<峤#�A���{��r-���j�,�<XU�C���Qm�]��}#Ӷ�\(�0&:�$�cy�Ȥx�-I����5NG��t�Wx�
��Z_��i���juB_�*���Hh������V��?CgУei���Ќ��O�>3�`��[�Me�=F(S� 2�)�]��)�����(�� Z_x�T�q	"W�y)���sH�%�xۊ�K	��H�����!J0B�5�#���i�4��A�؋�ć P8s���i���_ֈ��kr�*�\�&Ӏi&T^y�8�$��#"_UG� �[����g�m4���\� ��̇�	�|MJ�y#�2pO�����V|��ϸ^�u{��q���%�E��PS�8Q�ğ�'7��1��r�Ga�	�J�z^�la�?Bb����
'|�.�W��8����2�\�T�؝���
:F�ۅy�e	x��qT�8�~���{n2�IL|k%[P���&1�>(��NW����	K�ZA5N9����}���#m�uŘ�3+�/�K�'��ڤ��p��Z��I)���M�zqA�9޶
NQ���.d"����C���z��N�`X�����k������2��C�|`�~��|�r#��[�H7�8�����?/b-���ij<;π灋�_���������:�����f��@����L*�LRc�����XlxVHYEB     f9d     6c0��	�Un>M��ȸ=�?�;�8�.����E))7��q1�EYǏ!Z��21îW~D���dNK��L� ^-������+11�\�E������vL��Q��9u�=�H�����i�m5��y��㱪OY���|�/y���2
����P�?��4nq;Z����1�T�nj���f��*Ca;���+��p����.��o����l�4A'�W�*�m����-Ґfl5���Hx����|zQ����Q�5�&� p���s�>������̒X�I���Ņ�=)�!]��W������~	,������n!T`��/<��`#�+w�(��r�84�5�*S�*
$��Q���}��ϐG�F����f�0���~X���w|��wN,%T�%���N6*�
����ue.t4���2�$�D�sF!h����Ly�KF0��Q��4���@u�rg�w�U�&�|���6F��C�M#U���մ���_ �1��%_p�~����1I]b`C�ŝ.�`�Js/�.;#j��좎E|2f�����4���~@qAs?Q;3*u1Fr��	�Y��5�愴W��Y���8��S�XYׇڢ?��я�T��ZniRI��+��1p$�>�NT�����h����B��<�cN}0�+4�-LvA��&���i�U�|��c~Xt~��4� �M��r�{�N~F<��<�Tk?�ëX-/��0�d[�89�fe�Qc���l���n���9�����ެ��	dP�̧o4��B�i�f�d(����9%~b��\�8"���:��������q�Ӱ1�Ώ��y�f�SQ�CT͟Ќ�c���&�Xi�H�ޙ�1�H�@�59I�.{x�Ʉ�A��K���_j��5�F��v�N�Ԅ�L6��A�ǈ)i��Ձ�lU�%섎��lΙ�[x���~����A���5$�	�WS���<�R=V�4�����0,$f�yV!�M�M��s���2�6��[Uws۵��{�
?���V�9(Ū=���B~�ǃ^i�
h��ZwBq�ȷ$�SPN�7�/�3>u�-�ӯ�x�x���-�ܐlk�D���7��\
���P���a9
�+3m����G��1�`=�1�,ɍn�n6i{|��0Q���\L����� Ԅ����>A6~$Ч���-�Q�K�d��?��v�U����%��!���˗�a2�
\� ���m*`�
���OF(�ֿL�pQ%Hd�L�(��b���[%z�LcbUw/����n=T%�����B? �#o�h�bњ��O&���@�x].�;�.��A�hB(Z�LS�����J?��6G$�?v?��."n�cKH��KO��Ɇ�_7�kBG�Ơ�_/"I��|lP_[b���2�@�D?�pF|Q9f�屇�׭<�Wn��q�q1c�?g_�՜AYwb��?�J=�T�`I�"�|���b�q��q�5ףw�b y��Y(f�-��p��HO.�{"_��m���zI_�&��k�E�V�)�����5e����e�LEcW��ϥ��Z��`SF��":���q�W�&�J}���&�L�78;�N�,���r���-�;�JEH�j}lZ8U������R+ݵ o_#�jif��� ͔x؇'���\�y!�b�*G�Ȕ���Q!iA"�G`�% ?�5\�����PV�!���B�绡+�sD��rO�[�@MBICLq�zF��q�����>.��kϷ's3VOv��� �