XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��u�17���<���k{�<wU�iH!V��G���g+��ɖ��!4����3��)eB!A,S�L/8����qwAB�d�`!�~�w_J� ��mL���_�iӺk��   ��8+F�?,W����u��\�V=���,8(_�Ǽ�c)BTf�Q��+���&5�T�]�~~��z��d<�܅@S������=�����u�3I��]���#
z��tb�ʦD[�	��g8p��+s7>�aH���Ҷ�:��R��NG��6�)g�|k��l�Z��ƫ�i�|!�M���:�0����⓶eW�z����vU[�a��{K�k.�)���@&]|����jC�ݹ��^y��$�ԭH�
���ZG]�}��Wz��迋����������<]��$�Zc�~RMvv��m�j���>���Uն�M��(wOF�?G.VW70�^�!���/Y0�1�msz��p�r8S�WE����L�a��ɬ��� ���sPrd�]����)�Lv�·�d���3tV��,gi=�nw�Hw���L]�7:M&��|T��𲓧����.��	�����D��iѴ����n{��H��;�S �'#�KV3#-�o�H���֕�@ ����&�_�"���k��3��enH��S�����-�9��j��ҷ&��?+凄E��Ä��8,U����Ǔ��1~����;{�*�&5�����,b� 6�^&��?�����(�k�
�����XlxVHYEB    5866    1100^:G^��L�tԁ�em�LU�/�7;)6�>��S2�Y�Vg��C���ʗۛ�zz"pE�����v�8:r�����J�~�W\�'�5����J$�a��OB:�ͨϦN�e�-�SXw(����Q���!,�u��g��z;BYg�[I��Ys|�pi���.��(����g$OYz��[���r�3��2�z#!E�~ �D�Y$\��z|g�+{��m�ױ�Ƒ�͘�̐?�y�,�|��lg��Ve��8&���WF2ؼ����g���QH�6��e�y%N�� ��!�j��)�Xi��w�6��Y��N'�.8n� ��(�u���5tS~)!#��ov��4x/àLo��c/�M-U�U�n����k��P3$hc�����Y����Y�W�س,�r�j����܃f�I�=�y�爠C���l��%&�V�*ݘϻ�ԒV��-'���,���|�i/��ѐAY��?�����xzR��$ĸ�����c�Ɏ�{	#]q�m
߯;��3�f�tO�2m�Q];��R��Ě�=�K�y�T�XX>�]5����2�%CmE��!���R��"��U�}�V�F�:]/���L�w;t��;����}m�ǃ�$��w�℘j:l�#��?x�Q��YCA5�h!�H��G6q������R�3N��2]�t����}b]꜉-�qUٗ|H��2k�o�r�:@v�e�&�ά��5M*k�$�#�=�? �J���;���i7f�U�n4�2un+���=�3�܃4��aN�5�ݾ�q�kl�Z���nr�Jkȕ`啬6����h�+�Q��U������ފ'G����2�ں]{R����*)� �F(Y��%-�r���b��&RDeE/Ysrzu�6<$:5��;p~�� ��=�W׽?=�p�Ț��N���K�5�?$���	�w���KC��2�~l��'y,���j�:N#��>�EøpR�v �J?(y�#V��ibh���D�����˙4�s�p���q4'�h���5Ex����2�˨Y���a�4*��b���cv��ƞ��"Ȼ�[�Y�*����NR����(���)�"��F�B�kL����*���gr[�.��,�F�P�hA�l��n=�l��� f�.��v�r����'��9ث�ٸ�v�V�s�˖R8��98�	����
6��Cd�0;1�ؕ:��x�j�J_�VW�/�_l��^�(�F7��4���֡���k4n���� ��5�?�t�>�{�s �Q�+��O�z����)�'1��7������A*9����c
L栿	�* G�`_8^3@���m�_�l�7ϕ=�m7l)8���}���H 9@]�5@D��(�� ��Pk:��[�d�A{}�-������¬��pܺ4��+FiQ+��"��3 -��g�	��%�6S���5s���TCd�i7 ��<���ʦlg:=ʽ���1&&j�M�A7�xU��Iz�ggT����I�-����6�,,<�ڗ��X��9)~u��kC{i{��\<f�`i�1�w'���W-�'���7̜B��pz�Է ��n`��\�C��\.7a �=�C"r�;�9v�7cL⧢գ諘����ϒ�������,�X�d�Zv4}]n� ���K�RZ��1b8��K`s���?vډ�� ���R�@(��|�OwQ�A���	O
���+��\��h)����nB6�vP�sr�2��6q\������W��wF�z7z��!�ДǦ��Tb�$/������DT�%�t:}��'"2(�s�0>2M��7Z��4�YBYy�C�*Vt4o�ǡqڻ3B> �d���9ڝ˯�9Ş��#�V(���.�a_&���W�-�J�_Y?�U���+T�(`�h���Gƅ��9F�ر���t��F��*&5�,�v�J�:���^h�
�WX���z�h�:|۾���i>�$:8��>��x�����F��DX8n����<�`�F�D�臩�au���e_Cܕ �%cg��ͻP�?&��}\�_ݑB�C���k;�_�g�!U���+Vӛc��Z�$�YP·MQ�M4J ��K�r�ٍԙ��|����j���m�(�؉t�B=��ޚ�+����\�u��Eb��Ĺ
:�%:]�\�ֺ.帏~B�������2�:;H)�[sOB%i</�ca�DR�ӍG��D�'3��=9Հ�p{p ��l/(�	����u����7_3D��]���="kO�#�<�͔�z
�#8������O�{����K�K)H�v�&�$ _'e&��P�om��)'Bo�qb�J��k��4�v��x��ݹ�����ZNx�O�������4SU�GT�Fu�L�V����HY:�_<Qoc��ž�Z^T�ʈЪZϣ���g�!�#���������\���j�\mvO:�k���Љx�z`+�oBب I~(�12Z����p�B̲�?V\m�T;6a�;�vk 4g`Y�����Ҍ�#��-ɐ�D�F30,�y�o)�L'�y��Xl/���~K���-�_�	^.>/���kV0��?�$�.��a ��	�-���J����z��v���S`b72��
�CA:��F��p�K�ӊ��R'��4A)�aXMx&~��/�
�G@O`he����5��Ԗ��	�K�0^�߇9��n��y���o�Gtx#����QB���IG_F�ZN�l=lm�=�,��='�N	Z��M��00�c�X��q_��m��Sdv�_v�ݝQ��`͉�0�]�ƶ��s�E�]�2d%��ii#��x��֍ (C�l��v*&:E}Wyt��) �n;�kr�Q`{F�c��Zx�_q	E��qF��F��v�A��[q�p�W3������O�UO��/�mDJ�4������H��'�z�w�O�֌�H7a���U��|�5�톞@=3(��qAT?��O�i��=(MHƹ�t<���ӬJWǒ!
=(aQ1[Ѝ��}T�#	7���'J�m�<�P��1�doJBԄe�k���\T�0LJ[����h���'N�>�t�o��\=[g�s9H~�$��<��J/!�ȎATz|�g��<=��� �6���`3"�������=OF{�B�[6�{��1�M�>�DE�#�V;T0N��Ďi���6��k,��RM�j�RT���D�t�]�bӽ[�GP6����s�lw��]���������v����ox�4�O+��$*�C�������Qp�+��+O��1B���:��1ߥ�������6l]P#�g�PU�.�2̟��vʷPL���V��D/����#��A��}�1�N\?�B-Ԇݼ0F�.ʵ�zҡY�h͎̺���"zĬ�X5�?�wJ�^:��p�+<�_�;�s�Ǭ�*]����@�́U����/�x���
?���dnCZ�`����#=�li�X9��@Y��-�ˁ����^�l&��^�!���HѲ�x�;ִ� G�h�H}�E���� �R�=�y�-�h�<50A�h
;|l�)nNA��_��3�F$�2ʂ��FD�;Ǽ�a����'jPa�1)�eZT��&��z���;�i?�Y��3>@��v�nn<��-�%�{����A&��0G�	�o!iyV+�Y�������$mҷ�����.!>�{�;L�MV�Ďf=�.�N��_��VpSz������Q/w9V~�C���Q� �!{�+p��S6gȵ�移��]�|Uq(�|l(��[��������g���h��N�x�d�~ԯ}��ܨ�4�2�%qP#���f��9OL����p��Lhb	��.�e��R#Nb$	�`�y��`��cI�C���=o���n�#�����W���a
`�s�v+�7W���1�d:�O(Җ� #ʿ�x���ߓ>ȴ\6�U� ��?��F���)�p�cm���b",�f6��6�F7��/��?��;��H�c��< ƞ��d��rk�)T�8dy�y4���_��u�:u("�B����'
�4mN��#�ݖ��:��-�S��[��&��H��R�Ag&|v#rD��X�����y{ �2蟀������v���EFxY�3ʨ`�󞬅zQL*؊8�n<�n.��H{���xΏ��hx�Q1�5�� q��7���n��s��۰�9�!�EME>�Ã��Hcv����拙޾�@���Eڻ�� �pvd*Pn�ֿ���6�1�Z