XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����˳
���Q��̺��T�H�ADd5���E�y������ii��D��v!��47_x���"�;�����k�Q��4�|G����ix����6L/#�-Fô`���z�ȃ!O4P�l�=�H�`_�t���e�d8�<�.�A�f�HF����V��˂�0Uў%'Y.�nf���)���7Ny���ZQ�����o�_ft��X�}����z�����黣�x	u��D]�8�ĸ�Ztݯg��;O�Nn�t�a��Ǖ�>�o�\y�p����R󭝹���@e"i�9hhIz{V"�;;�%�|�G��d���E8F��:�z�^��A�G�l�Թ�����=��6D��K}k~�-`a."s��R#=v�D��J�憀���}���I�ٷ��#�^����Z�K��`t/| @�����v��,�5�K�+3��
�j>W�AV��}\Q�v���e^|��;��ZC{mY����#G��</�6h	�~M��q�D����Z����ii�g�H��@�^�i�\w��P
jۅ���"��~�Û�x�CV�	k̡=kH �z��4�%q�H��O:C��q��c�JJ@�rx2Տ���K�G2Gx.���8\O2������+`�]�d~X�cu�����r�f`�����4�!l� ��s8�*��u�r�;?�T���)� ��e�pv�,��[,�c�LQ���@�vu�PkL-��h]d? �LV�kY+A��J͚��$1$Pk_���U���>��XlxVHYEB    3c24     fe0��}�D
�q�7��4�|�ק�>{��2g&�Dg
G�^��Q��E-xc2͓	7"����.7�T`�U= ^��������7˯N�$o,@����ؿG7ޙ=%/6� T	U��I"� R�I�I��΂rv�0i=6���k�þ��Y���>�B��c���<��᰼��0,�H_{�!��Li���dN\��f�v|�I�"_��������e6�p� o��4d��W'�<�=����{�c�<�g4�;e%��ܺ�.� Q��Q9�˘� ���iCCJa��'����L����&�y��nf��ja��:����J����'����U�/1�����{�#��Z�7�K�Ưb)'�����3����0x1�𱿈�Z��D1��98O��*��Y��} ���8������u�-� �Q)3U�^S
}doKK���"��`bC�X#�ү]����q��yl���B�����E����.[�,�a0���~Q=�.!FV"�=('Q��h� ̆��\�yy�Ev�;�.!��b{���)�_��ۦt?y9o���^Emj�u�׸7k�&���hI��Fȣ� QL���Hj,�j  ⹈^I�'�q�I��<9��uLdd�����qCG�m~�w#����vϹ�.���e,c�O����y{��8�\�sW:Zt���Ey�3���	��|�Cw�v�i~����ħ)�� ��I�S�_�L�;��q�
�2��16�&�z��{�U}F&Cd��U��v#��K\�<dʧ�qŝ݃�t�Po��n�w"$x�Gl9Ι/a{[벜��/nP[�\#{��:r��ߐx����\8Wƽ=���j��I܉�6�13:S�J�=>&qS����b@���[����F�A����g�h���\;���w��.�vw�����j?k��-����b�y�>�W�T
x㣚<@���E����G� �[ɞb��C�ׂ�Q�h�M]!W�q��;"I,�<{C4��#��g��
c�it}�#ݦ�A/^��X�>��QW�_	'��3����4�z��a��>H6U���8`z��"��������G���a,��Qn�Up�B M��,��K"�5F�_?d�!�?4r�a�:��CU��� Χ��V�K�&���9Mg�S����:��M�?�=G(<�=C�l"�X>��L��_�Q(N;_t S��ۈ�q�h�A��6C�U�ܛ�|�!Ӱ&T"��3>����PW�3B"�����`ow(S�d|X�R�X6��<�F�u��Y�Y��Ia��5�k8�+��Ej̓�-j����5�컄�bt]X�X��U5]7��M@js�+C�|\B�k]�V���c'~����Q��Rp�f	|���+�pu�9����-��, %��>�rB)���^g�����&�ח�x*�q��Y1������7�o��jEl�a���*S{�c��J~��ǒXO1�ӵN󈘳�
�cW�B���
�9UW��f!K���8�\�EL<�����U�9���(Dj}h?���4����"�`��XOGQ�V��ԍ���ѹ���&�a��K^{X4Sh<GY�@��x�W� ҅L�;�8x���T��J�8Ã�����5��?���FOiE��BKJh�.�!J~A� �9#Z�t�̣��PH�߯�8���=�Eb�5l�+�a���Cd�+	c�%�cf��&�M�و+���[ϧ�m ֆ�ѷ��5=aĘX$R5�����"������7�H��y!S�@D���o��p��H(�P�Gz۩؉r�8��p�s�|�#�������8�Θ���� �( *�
)5�7g�|5�^>r��5��V�#:P�]�* )��:>�q����f�����b�s�%=������WG0×��ν��>,���u��%�ȷ�I��ĕ=��Z�:���Cy"&0W��5�`�22�.gXUGN+x
g��$����[�6�>�Bp��V�6]��(Jr/
�zV�O�d�D:���*.�Z�a�)��f�TܼR�"M�2�6���u��3r<�eV�ъ��Rnu�������S�Zқ:��r*��%2�:ͦ#������N濅/Z��y�#�hv2��&>�y���B�Z�UC������V8���Т���<=���5�'X�8�����o\����	�P�<������i);�Ʉ����Z����g���v[�%~Y�OO��F�k+�h��d�? L+�m�aV��Y��,G�Ы�P|0���	BĜX�L����A���3�
���b>j9�x��"���F*[�*6Ii&�pп�����&;,�Z8$�y�5�.����|��c�n	f:��&��n����u�qb�Oە����+O�\f�)Mwu�dǃ�1�i��/��~�m$���T�XK֢ݾor��T�v���Sc���`f�L0њk��a ��i�~�_d�~�' F���l�E��ʍt�\�wS �b0s�̫�{�2zy �>�<��
����m���-�!����"Z8*#�ʎУXkMME�b"��N��ii�����1Ǣ\�i��Sd�(��d��X�{�������g{I�d�]YP�2�m�������Uc�Y{�b$��)�2�L��N�Lp:힂���nE��D@���U�qq�c�#���HQq2�qpڏQ7+�JhR�b;�^�&Gl.���I�	����=
"J��?T8n�\�l��KIX�YA� I�yO�k�0.f)��b)k^�V��c7E���'r��]["u��f��_k�:�My�[Co&����	��(u�[b��/HH���Za�����5���n%��I\$���_�����_�p�m̳φpo>?yN�Z;Cf���m��\�n��ѥz��e�� ]g��90���f?�^�bߩV�)�j��'�ц����4�f���
�_���HJf�*,mZr�oο+�6R�TS� u0�=�X5+�����b����ctx�k1�i@�:�kfC�`PRJ�r"�F=�F�E�t�s # ؊��fXe� ~�+H���K�����0?hM�^��]��T��6� W�I�|�EI�V�D˾LHP�~����+�H�(�Z���c����;:q(�'(���?ٌ�.�r�K�M��#W����d{������oߊet���4���p=�����}9^t����aǉ�Iƈ������4ʞ6��Lz܀��J[���	D�%l�&�ڪ3��欤����iQ���ک��D��1�b8�����۶W��� p�6��N;o���Cpl��P9s\;��U
	yH��R/I(ث|��A���\�$�!;�λ{_�H da���(�N��~$J�x L��[��@��K����&	��(�٘>&Z-|��f�Q T��&e_&�0�
��Mڹ�΢^�o\�;b�4��[�i��=�~����Y���X�e��\��Ͳ@Ϊ�v�O�Џ?�<��d�J����!:p"��~h�{ ���l�ϻb���n%@�<�*`�ܓd��0/čw	�s��.lzc ��T�5���R`�<��}7�N�=�4��"���ҳ�]��鞍���6rzA����[�`��d|3D���l<�)I��[�"��fT	���^��B-�o���U��m\(��{���b��X�6�ci��$�h���E���}O3�)0��S9���IG�c!�o9/e_�4�(d����s7�?��=�:��2��mB�'đ��~��9�o�G��O�՗K:��lQ�� ��2��B���Z~m���0'~��Z=���;�dR����H6֢4��>7��K��Y��Y@L%���*du�I+�D�΄L���"��z�n��nU���s��H4��	���-�vzR>J٭|�N�n+�]���)f�R4����|����T���m*��	�ǡ�/	S�{I����|�x�����Ɓjy�<�������,L*�h&yI�2k�z��ӷ�|���K.�,�xi�Ñ��u�I�(f��g��v-