XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������
�˵����m�+v"�B�JI�.�ν�~�n�����ؐZY�,�|y/�O?K/8��V���z��>��8��`^���pP�׶Nu����w��EsQw����,a����r��?Ӈ
�+���1N�몡,�/\�,��XQ>��/+m(3)Zc�4�$��fp�>l����{Ѡ�naLP	��x��f���]�$J�VX�ױ��}L���|�=����d��T����5Ђ@��,,3w۝e.��ْ3�0Ǵ�A7R�Q�T�C�g��?����z��v!a��@��o�}�{w��l�/�VQ�ZT����$�B���!qڵ�b!0=��>�E%���a��	�{�x��!T� ��di��G�K�F���T�q��|d>����f"�gƍ�[�ouY�(�w���J�ݓ`i�Ij5L�"[NW�ѭ���T�U5��"�������0m�̞0��s 9Y��9���D3^�:���\��\��JJ8���>"p֞�,Lt��}��4`d7������o�풅��|T��#F�bV��x>!���?�_��ThY����>�\h& n�F��)i< ����F�RS������-��`�RY��p�-^��ȵzÃ�����nF<�r�l���N3���Rbi� >O�>� 9�RM~�'@Vim"f� ě����K-���W/�d���x����J�pί�f�����7�b��	͘��8e�o)bEѪ��=����YH�@��Hf��P|�&jpY{�XlxVHYEB    dd8f    2160�&��<מj��&gߨL�vA�����jc`	���.���e�l6�KX����/��d���ͱ�%N�B���`<+��F�sM���YX�����B
��7����Ѷ!k�eg����8�$�Hol��v��7��6��Ȼ� V�1O���� �[���V�	5��ϩi ��$��5�XKCP����xÊ�Ev$� ���k4�&i&�s0� ��m��0Q2_�f�:A�58���L��[�l�����t���wCT,a���
�S�?#jA���-���1���igƷ��|� ���ӎ�Ͽ{eT�J����+7������w�ΘH㈔�ͱ�"l�8�x�A���;S~����]��D��*���OFF�NF��aY�l�2�+�����i�4����
�iE�5/٤�z:p�+Թ�HF�K���M�sL���UOj�-��g������c|(���d��H�t�,���7��/�~X�aV/��jn�2{T���Q�MI�<oV_�L��YZ�_%�����B���s�v�HJ�/ �O���tzj�ۻ���M�������c	�+�����0�b�m��b�P9��0��'������Ύ�_�6G��2ʄ������ �.���{n��St|G��_�\M�e����0��-O�q6$ie����4gD@p!�j��>���Ch�«&��BrFސ��We������~�>�%#'r�nT��f��#x"�p�3;f���%&3k�J�l�1�3v���H8�O��63Y�����`��R]�� fI,�(Bf���
'Ǝ��T��h�z}�7v�i�Z]��x�����h�U��+��/\yK�f� c3�a��$n�\�O�w�,��`����
�2G*C�ŏ��^@���I�W	���g�����j�A���I�'*��:T������"� ��TM��~S�gV��y�vW��!�:���GY�x���*6�#_�Q�7��oL�aX��۰�#��2��T�����4��������"êpq7�T���v��_@<�pD��}�͚��2/b���:d�^`��xՃ�2�I���8�s�̰��7�X�C��%�0�֟2��Ƀ����Yw��>D�\�U�T(W�C�%q��_�d���< �<�E�e��X��J04�ލ�ym9lu�[�=�ԱTC��b�{ԴװF���-9���IbW�5�c�&ND#��)��MY��I��`�������� �r�Y;~e.o2A���5P�d�.�E�����+�{�wiO� �(�������<G�V��ͻjY��>�U_���a�$m�2��nq-gm홊�&kE��1q�Ko,`�EX\�,u=~M޵�p�����/��Y�)G�}��f�>gP
�T ��&����e��#�i�)���־�9��͜���*RY�߿��qF�y����8��(�HZ_h��O������"6�����Y��6��8F�.!�n��T]a�LJ7�h����)��$�����@���p\��^�DF֎��ϫ������F#�@�0݃��-*��bj_�%��-r�/��fsA��m#O�T�,j��N![8䆤1�,W�R��������Eۣ!�5��-��ħш�]��2`Z1k�M���U3��SVpv����_bu�r�[�)b��r3�P���e�}&�s�:�����R����&���1_����Jh��X "�R`�"�.ّ��˒vĹ�[��W�-�ǂ�b��˃��r�~>�����m.<:���h݌P>W
mh^�-�bF��+?�y���hR���12���=�'xj}ܼ�|�{8M�U�cHg�5[*u�2n���Va;������51�RS�1�3�ޒL�;�;4b��Ҕ߬�R~��W�|�%��ʻ�oF���� ����D\-����G^QU�>�����~7MO�i�b��?��Hj��KȘ��%t�?O�<�j2/�&HD�������S�����H!����7B��Ѿ)6	p��)Hg�{�x�=1)&Bs��1��,&,D����b�f��?9�fTڝ�;9N�Yn��G߱���`��c�Ó:#/��G���Oʔ��S��CF�!�����E�q1���g-j�([���PTG�|���q��f��`�UIT���l%������T�wS�|�����Z�@eb��U���@�jS^9Z��XL�z*�<��/��پv��7Ej3R�Ć��� U��`���/8^�C$�x@�f��1<�����'k(k:=��c�$�El�,�v�a�S1=��XQ?�p�5*�pT~mM����	��F�Z	']�]�׺�N�]�
�����o��1���$���^|S���o�.dW��w�Qg�]�b'ދ��8���|�7��ƙ#)��qʖ�d��( '2HA��G�r�o(�<�q���漷����>Zx���j) 
���[������V�5�%Ӝa"6��~�R��!��ȥ��;�np�9��h���<��F5�p��܋�N�p�-�b�V�Ō�|�2>����(���M1�bI�!��9I��ޝ0�?��Ȓ�B����fn���b.jGU�1��1;ɂ#O���g�46�j@P��j��@�؆:p�)X�'�j�b�Yٙt������_pV  P�k_��EVJ0Q� ��!	�76�^�zO �*1��y!����Gh��~ݱS���Ne�Jx e~�9�V�4��������Q}=��9 e���9p��}���h{���4�]��ǣ��I����� ��`� �!�vg��w���[�Ys�V\���=��r�,:�}�;�0&$��r˰���<J;w�NM�}j��[�y��#�4�\EpYH[�- �A:Q�W�#>3�=R��(f��G����}Y���p�8��5&8���w���<�G~o�o�c{���2ݲ!$��ҠT��QӗX<��MdqX�VyU��892��x�*?Q��-�9	݃X������yo>�7B�����
}{1�� 1��ֻ鱘`��K�<Z�jR=�&�g��>���L���T����k�Ld>���K��K��B�($�>*�%��n �.�٧:�q6�Y�~�;�)����;{ϑ�k��7$鹠��}a{����L`q<��q��Y�Ϧ��U]Β%4�w*V~�>�~*����$���y��6�y1B���V��
�{�d�ǰn�H�;����2�9���12pz`Pf��S���l	�c�z��[����e�����;	��.`2{RX���-u��0�g��+_S¾����u�eȡDG��4����d]*������B���������k�����ܰ.H�?��ߎ�鰷Ҭ�yZA8���-J�H�sSГ�@�������C��d]�D����i1��V�`4���ݭ`�\>�NE��e�Ȃu��@5 M�j�?�x���^���r�l]D�y��e�Ty2ĳ���؛��)C)I	�D����V92��4��8�����ڡ�2�$Ex",�;< ��H{�N��S|���nz��q�p�&�����tð��S @�m[�$#d>IH��Ny�	�"{����e�
���E��y�F�1'mm�5��!��t�(f�s-���&pn��^��˄$! �y�=�*ӭ˓U���ίr��,�o�t�����o	98h�X�5�@��sX놚P���ıok�����J2	Z���i�c+d��OT�47�����k�˃�y�:�b�jKCd� m:�wޢf�V67��m�^8�0�ډ�&Ԋj"n��\��)7c�4�5��_M�1�7)� Ǝn��ݼr�?:�L;�������G(��o�$%�E�YV��I���ԛsv�o\E��6���wH/��i �	���)��ވ	�O��]B���.�Q<��6N)�<��wm��ڊ��'e�&M���������B�Ԋ���ƀ�8����9����9]ha�}��<j�Y�2���F<���$eV��q+FM�OCO��nAcjL�����Ub���u$�)����Rh���O�x��w.�&/'i/��h�x�<����@�`�;�.}�W�*c7���xa���� �0'�T�:&�45��q�Nn���(���u���Ni	�����Ú�D.E�jb;=8gN]���C06�f�l�9���{ �J�(J�����zG�e7+*�2�S�9v�ʹ�����w�Y�p����o�e<_���������8��w�:�:��t\(r��m���Oo@G	�|{�eJ?�W�#�w2p1��L{��#,u�N3�򴋎�x@�!���0Ѵ�=$"5O�ȵ^�mG���i�Zx�_��C�{l��r��`��rβ�����=��^vF6
!��h���������Q�������!i���[�;P���*�[xތ�O�X�H��{U����؟xF�Λ	���~����:{笀�u�҆)	����S��c�U��@\.��>a��f�NeA�~��E�sG��o'�ٞ�c*�y���N?����h��_A	nh�X����А�ek��+�	L��g�4<-U��O�I�u��>�L�IV�,B�iQ��{�6�z_["�m{�I�Q:X�����{��	�❆z饐��T�1�ViRU�Wl6{ўn�
t����5ӚK��x�z���w��!33�4QЈ���y���DS��8�D�Qe��ԭ�A>w��������rM]��ؤ|m]+]g�`�~��: /s�^��in���[���3F��'�S Nqe�vh��c�?/����H.]��3�V���sE����&�p3j�ıҗ� ��(���gI�|؂�Ь��0�B��pF;O��	�F��{dP�I#��C�F��� 4<+h���'���<%�N7��Oi?KK���Գ��{X}�M�{χr�6�Cr��$��~��@�C�0�?�}n���u�h���nn�!���̓*E��)�멡m�-��d9uV�w?��֣PA�"�)i�T�z��SH�68tA[�b��bS��O����SRK�	"cmo�k(I�JD���l$�#q`�75�RF�BW4#�l���nR'���ߵ��A:��0��dZBr�?�)o7�:��t��秅�2^�/�F��"�U��[TFqE=/8&�e����I$L%	����^)pF�Z�S �r�ߓ��
g{�� ���K����2��T2���Z��l�J�6v��J�m�o|���Xx�*;�+h���F��"�;�ۧ6�s-.J5��c�(��d��N�o�:�q�<lV��٩������=.��₾?��r-�=8�f�k���Q?�@9:�������:�Q~@W
"�k^$_	��U�<Jԇ3�4%jަm|t7'n�=Ws�����B�{�^�;���3�f�j�KI3G���(N�G�x2�
ῐ�5�x#���ˌ�@����<��A�kt�>x��8�t�\��< 8��T}�GQ|h#(+�"��8:��bN�D']�������ؖy �#��$�v:��9���s�\�r�B������~y�
�J�M4��b��8�8��gۣNlYP�l*�S�"���%�T�؏�>�Wo�M&-��QW/°h'Ϝ�H��op�j6�=bh]*t��������5����W�E�x_�{Ȅ��Oڔd�0����k�9��x.n5?^�ʠA)�E�.}�ޓ�<�0��)��Χ�=��/R�����#�/�J�K��e�#�,�d*���%H�W=��!Y�2��z�nE���q�R��!Mdg��sTx����	a� �J��0d���x�?G�Yp�Q	�L,���qv�_̑_�����;�#(���e����C�h$�1��KPG!�"�����e�Ѻ�|C�T��]�����.�P}Ɓd &qE���#�|������Ď�|R%:'#�\�ɜ�o����Y�0�Y�a&I>��'�2�@���گ�������O�^�H׎.��=4��y|���)y��L)���&��[�Rpi��6�	p|X��^��"e�:;P�n��������m�����4 ����&�7��� w���ۑ��> ��}��^�#�8G$ԘX<�����Y�NCL�b�{>���B�B*�m�K�zz\̧����?���e�"� �SĢ������{4�50����.�w�����1=@��f��K��/ҍ�L48����iDF����N;e�7�j���YI���#κ�~a�3�a��Q�e��wPyo?�����@�q�Y�C2����}]V����0v���۰+8���$�M�_�0�.}{׬�2�R�Z�"M�TB�9�=;^�.4�喭N~�(-�_���/�]8����J~��N]���=�0�DӤ�G�-^�!�&���w���d��++����c>���؏��(T����v6�I��m9�&�1��.����L�p���Y�v|�<����"���cf�
�0�dt#�_h`R��AC�Ū�m����,���ݳ}Q�@M���-�6bg#Y̯Jy���e�7 "�4�#�{J��]Ip� /��( ��|gTo\�7�p��i>�������}�(�C*��y��`[cq�����C���m����JG�FLe�/F��ɖ��*Aq�H��yJI����-a��e���D���3H��t��-M�|��yǞf��YE�)��W����4�z�a���>�a2�0c]Vڒ��
"�Pjr�<��2ȟ7!�Jhe�ؔ���������ּni�tR���z(�<�؇��+U�p�D��JԳ��fIˬ��u��"��Yu�llQ<�^x�����x;�Nn�8�K?.�Oq�]$WV��K�vVӆ��=F�n�)0���u	��/S�i���ޥHG;0���E_]P�d_)��~�z%�i��1ݺ�<�4f��[��mm?�M};�v�
�����v���������㬅qJ��!p�%�B����^�q�~o2څI�6z�Չ� "C�IPl7�emH����5qb�R%1�[�S��Em>�Q��o�^aU�x[���-�<ڥŭnxA:�q�2�����������R`��'�ag���VV��of�qI�5eV!:!�>E��jt��'�{��01��M<K�B�k0�5-�HS�G̹�<����*�������>g�t �%1�tH=����:a�G�Ӿg�ЎZ��W!�Y���ct��l`:ha<"gc���˖��{1�:ݲCC_tr�0�Y�R�%��~�0ym]��+�%����w'�JTH��K��i�����%�a��f�͜��D�S�Ë%�ϊwt[Ch2��pI�~w��tݻџ��ϸ$5k�5x絕�y��Ԏ����g؄�������fF=!�0�`Nx�ii��SU�ŋ�$(Pi��C�޲8l���8Z+�(�NF�}��#n�{n/����<ܨ�s
�.��d �D�Gi�-!-.l�N�6wbv3h8����Q~�CHʾ(e[��^O�a}�����Е����@��il�S(Α��t\/i5���g�9Y�0��Uڸ���\H)I���F��3c����"nZ����OH:з�Alf�'�qA��Ph_��Z�y����<��FȔ1q�A���0a$s�'��=k00»H����՘���[���
��-%��:�cT]mH���C�����K�5G�Q���|��1���ĺ���8+w��xfJ_��V�1�!��vP<��:�.e�̞w[&6�ᡲM�o��'ʔuu[$�����r2��eݠ�*8��H=W
�<:�1j�qܷu�U��t��܁Ϥ�'쌚2@��nO=�} �K�Z����t�ODE��	+cg�E4�9�;��<įV��xea�]�1.m<ՙ���~��|Z8萬� ��^ds#סBH���ޤ͐i��B?�z}�,�Q����:��uq�c�=#���%x����5[Ow��r�x/��׼���͛�F�MȂ-�ruA+
��Xk�E:G��["nt�˾2�+�]�0',�ʮ��_Qϔ�w ��Ґ��-Ԍ�n�q�Q|I�`_������S��gB����M�tTo�����>0=��HnMgic�W����Z��l��A��bX�h�b��VXd��Ϗ/�ٯ�Z�EwtVWޠ24ѝf���0��}��L%bۡF�/��ƙ�ϯj�L>�B����"��ҞR�,�{Aͼ�5d�;��I�`Xa O�-��??���i`f�-I��$(�YKH����e.����S{A�In3b�{��q�z�y<rʥ��~��1�;g��|B��"{i���Q�vAT+3��}x?�G�"�6���8�2��{��*���=Mm6�8�/���t�*��rn��4(~8�q�F6����<ޗ�j�7ޗr�