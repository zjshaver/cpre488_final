XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����[�e�e�ီ9:�t��*G������!�H�~"e�:����$=휐�5�$6+R�Hj�?�=w�2�y�eƴ���ebgN�V�@�F�J��<?m#��-5W���\�L��h��^��H{�5;��
7�B��h"}�R	�eǕ4$Yňp�%ӽ��)�ઽ�����ֽ�ĵBJm�ȩ���ݟ�����{���c�����x�hd�)�Ls=����qѭ8�ȠV�Ǎ&���r,'����<G�D��&�)���*V��#R�4�m�"#�Fh��!+]��<_��?��=q<�.�J������5qk�6&���"?Z�RQp^�JzrEc����S|��+i���W  ��e�møZ~��Ŧ]�)�T���q [ǭ�#px�W�nv�-/�~ڽ���3Zm��A��g�Q�"����$���"/@SAp<��h�D���b�Wǃ�$wt	�lo�{6��$ VY���;r܋wLL�j,�h��To���1IĢ�"�مw\�~g�@�>�I s=TӺ�%������'`1�e`y�eq����E3!R��i8���d�\��m��t�ƀݝYQ��:dtl����<�4�>�_��Y��j��cS��r<@�K5�4c��Y_ }z"�d*S�}1U��s�m&@�5.�S/Hw7z���1�4�����.�B���V����ZN��c��I�
|M��H Ro��w2&�3m|r(����AƯ��#�K����DiO>aA�WЭ����_����v~�XlxVHYEB    4052    10f0k����ILpb+���*>CE�)ǉ�ڛvq��ᅧ8l{���TuiU�Gm[����P���MOӐ�����X�����g4�o�#|���!o$^Y1�k0'lP�%��R.�Q��_N~����8۱���9��KaG�_�Ye��b��Y���zSQ�2��w�v'?�qGR��VV��
����wM�o�����CW�����LϿ!��9N�ý����tU��L6��΄�d�}眿����1�ĘB���X���Ӻ����,�K��i�/�=�6-}�"�����C`���}=E�?�TM�i!�k�Jo�I ���N�ĩ��
!��X�l�Ш���o%��B��$�
æQ5��PjG������=���f�^��b{f#f�Y�NUX�%�k|�i�����68���oL�9�ܻsyգ��5U��l#���Ht&��zuA(�'�J�>�-�@D(U�����+.Ȑޅ5���4ʤJ�D:�zG���A ���t��(c��]����TU��)Qc4�`���M1�f�@�8���ަ�Lܝ7�4����v\1�)jfuہ&Sl��H�{��oO��N��<��x��z�������!	I;�ټ�x��c*�;,6<�<�{��+�qE�B�ú�t)rb_5���te�I&�[x��;	Oc�~B�
��JG����#%��?pJ=*��#�Iv��:�e�r��7R�^��7HҾH3m�7�Ү|TG+
��[B���Uh�7z��K�ZRp� |�z�!s�D���CwS4�� ���>AU�p��&��|������+�_cc)�%kg9��E��!1,�< %��m5��Uczq����s]�5�@�IxP(�����ή�]���*��o�_5���V�] �����2�B��z*��~R���a�_�o����|	#��#���/�^�Qח�]���
=��yp�5,m��YwF�1�CB`�G�u�����ܖxI4g����X�^�D*�:������%�V_��i�^�XU��O4%�y���?)�S¬�r��'�b�@ve��|B����Y��GӓJ*��l��e�ϱ��i�ZY������٠6 ��SH}�� D��;�?2SW8v�Ǐ�٧(f������_����"��B�.���;�k��Wv�I�a����k ��&�/ɴ��լ1a)��ɝ���\��M��D�-�gm�Ik����k� ���O��Ȩ�*�kE&�������fCyރ��wݏ����+�{80<�%@.:ģ�0-��a*��Ԙ[�$t"L3w��y�Q/u�6���v^T�d6!��ެv�#�Y��D�w�\O�[*{Hz=Ns�X��?��5��	���݅��1��{�,'���ڜ	a�f���Y��Q�m���7lF�[>�.6c���G<%IY��M�<La{�e`���!��|�a�����W9�p�O����eyE$�Ryj$o�:ބ�*�;vW��1λ���o��T��Nq���1�Q�2�v'������?�&�g-Yu;����Ϸ�a?
����?4%�a_U�ѐr]��^�����Z귍єG��}�C���x1��
�����=�8CڶBRΠ,��D����?*�lm�l�U>�B�h$�>��'�y���+	��F}�\Ou^�"�5�J&�G5��)�G��:�l̈	В?k��@�k�H��e
��T����ήe���ԓ=7{gZ2tX#�1�M�@�5��ش��.N�X��m��:��g��Q���"�~�	a�]B��7��xῂKё�*�~��U���=$3dk�޹ܸ�RS+Q���/��r�7���@��:�!���ޱ��N�v�'3%��['�����ޝȷN�)�v(`=��"�m�ph���֪�N��L��xt)E���۱��}����c*�
��O���ɓ�?��o}��\�S_��
�٩c�=闚�_5�`�v�I�g�� �Ň( 	E�[݅%��2���*�������2�f/����;&��⣽��+ﰄ���6���#!%W�-SR�rdʤ�yGjQ7��Q�0��ڧ��<>�f�
��}��ɦ���x���.D1ơ�����LF+�=�9o��"��*��7�>~%�"�]���!۫֍c��Qږ̍/���04P��߯���?�,
���=l	��#���1��������º�2s�Ӌ�9��)��2�j��@�������右6���v�&Ļ���i=�:m"*�����o�V�&�J�R�6=x��Zvu�}�@ (\�T੶-k�z�jw�@<�a�*�#�A.�?�B��+Bź��D03H��ɢ@���8zZg��ʯJ�XP/e�l�)�;���!�����K�Z<����w��Mo렲��,h���;X���c5R*N%�Mb4th�0��-3}�5G>(S��4�����#�0m�����k���#���o+����)�	q{��`]���2cK�De�/��;���~g��M��Σ�� r�����$���~�����#����X����-��ef���v����wm\������l�(��AD�f�F
����ice1!M�A�H�§�'��s���>wn�O��64P����>���8K�RA/�W�k�kWT�r��T���"��l0x?]�����n�/���)~��I_"A?�X�촊t��ݠ�R��[+=�Vs�c�Y�L�L�+���`��}�����.����<{[r�O�-��l����C��?]�쀯>Z�b8�%���8 `,���L
��
5x�eW� ���I\���;*�L�6G�Q~�^���1�!>
���%ީ�վ�����Tl$��X7R�;b;t����ؕ�,�h�����T2M��F��N���:g·V�K�_�W����ċ<L���G|dϥʇ/��@����Dp(M(���TP�)�0���P��*m�͏��'tzX�� w���.���1�w�XH/0x��р�(���3��O>W�N�d2+̨�D��tq	N͵�cK��ڕ�.NYt���{�V:������������+����~�W����]�0�%BS;�a�C��&ห�H	��<�N��ZJ��e��uC��}��W3�)�0Ly����\��bQOJY2y8Q&������l�"c�N	�Y�`���>��5�)�!v�lz����B�1r�� �t"���2"]sR�}>����6 �Aܣa=��3�g�`,�Џ0y�m6�X�LK��?R*U��!2��(��z�(�+�Y�}ܼWy�~	�#� ;j �����KL�;��Չ���l��0�C�Rpu-&����F��7&z�w�J�'�=�]$�5;��ǟ�A'	���Ҫg�[�����~�(����ˠ��V��Ū(l������)!"?���;���ܥ��%��rV�������8���S�)�p`F�/�9���7��Ɏ�2g��}؂��KS�V��$	䕘K>�$l}���|�@n�9�X��o�9e\#k_��wJy�(4T�0x���#Tć����2�3 �L��.]�=������ˆX#�߹_	8���#�|U>��5v��>O.�PJB��K�����i���r�@?��5�h����Dč�0yV���f���%A�*��aa�y�c�U�&t�MH�IW�3�J��'��O�I���w}I�uf&`��J�Ca���f:�t�9�JK���F����漡�#k���kZ����H������w��`�) ��ç�ֻ k�����0�"΀�����
�!�z�D������&�h�$�P{>:�.Cbݪ7H"]����}� ��)�z��'��C��p�q�b���9B!��|�Ǧn��w�U���j�|~���e|�R���\y��W�ə��+��Ϝ?�A׾�)mJ��q�z;�[�=��H�}�48oX�5��:���!E���[��n���88b�eU�Q�"n����(?v����k��(�ʡzwu��c�\*�/L�C`J$x�L�b?-�"���w�H+&���:��S�X����Oz����u�H�(H&������h3��xqv�t��8�  $s��%��װ}�����2�w�����I���=-�'�=����k�,�xg���t�É*��h1v��}��l�ߖ��3e��㝴0��	'�1l����]��;�1^���o5a�9��=cnf���ѓ�D
$�I&��%�B�)fŁTK���ǚ�N�����@x����Hz�h��