XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����(�I�'����F/h��/�ӭ@M�}�\��E���x�C0�D�"D8(�1q�TO���N9g��G>���ڳ
�*
�UY��}��ؠ]Rl h��H����C�@��|ߐ��m�ef�b<�����m����g�a>�M�kNS�
�y2Fx�p0�Q�ǮK�To ��qS��(Ъ:B]�0�����Z=�=N\=a�h91�Ԅsʻ������	�嬆��n�U�6����.����U�"�^%�t%�Z;�`��>S�]�3�sJ���\GBʌf�佭�� W�2�����)��QDxK]���B���ыb��ۼ���^O���$PQ�E1�rN�r~�������������c��]xM�-��*���<8��F��_C�.�Fz�uc�೮�scw�
s程TFT�-&�hM8rM��!�����{���H�<���
�h�?OD:���|9G��|��t�#�dx%�����ݒe��?�����`�z���P"��L��Z�I�w�3�i7�ƽe�����\�9[�z�Ny	w��D��L�el��bHg2&6h
Y�r��8��೭v�쫘4D�c��Mx�:4�؆�-�=<�F�o��'8�,%�=���G�+�4"$Q����% ʵ�/u�c�L�yR�����a�Z&���c7�a
�I�I�Ce)�%F���[���'~�����u��Kg�ǎ�~W�*�����(^u&��˖�'�k�g���>�gP}��(����p�-�~Ju��XXlxVHYEB    95d3    18d0�>vt=ux��Ě�Ίz�!���@��G>��Q�<��W
�o�[P�v�uA�8�� �������n�.�in?�����hf	#���2Y)s�E����E����?:��~ ��5n�gՏ��l�nY|#�*�=��y'ҵ���%V��D���V�T��g���P��xW��z�m�s��� �yؘ��赶)@k!����mLP�0�*�]�����9��!G0q�����'���A���L�.�w�* }�;�خ�$�����f�#�5���@c�m)�`�7�K���u[ٽn�7G~[ϔ����
d EV��%�90�	nl0�OI�dqO�+��$+�@��4{�r&\�å����8����ݑ�j9���Z����]��Q^�%�ֵ�&������d/�׹s8�Y
��P&w��HY(�_N' � K�}ZHv�a���f �����6+�rK�t��b���?\���-]����?�d6��g���)f��Ǩv�!6�w9�.H��?�!&���`QS�y5�<9L[y�?����t�K���mFWb��ߠ��DU�BWT����r� ���Y��4�%��lD�Vx� QL�`��ZA�<��o�?Q�t$�[�[�޻��KB��rE����ɛ ���ˁ��#r����$�_6V��j�]1�	�M�\l�Z�����(�wQ�*�N��MsGs���C��VP&*����ٖP��1�!w�խ���>	���ɡ+��?z��5`2Cġ��<��(G� ��C#[����+]Ȏ�q;؏�������ӎ*L�>+�<=�F��)f��i�r��K-	�Z�
 0"":��ɳ��
A8�wqM��G!
�IR�gC��������z����v�M��0��4��r���5кH�@~�kD���9�HJG��w��a�x�ѓ���~��Z �|v��/�ǯ���$�ThYC8ސؘ�#B�#�ӫ�s1M�I�f���,y�D��s��s�H"�Nv������\�T8�K�����Ps�D+7�����5�L�4{d\4�`�ds�
�b�3���ԉT�������"��ex�"��39}>�"ZQ#!SK�v�����C�k���*u��S��N���02�t�^,I��`�,��k�X{E�¨j��:�l6x��mU���g��߅�:�������lD�'^�36�3~1�>�D!�㝋��M��jWL����2�����cfN��fxA� ͓
�\oS�w�!�F��;K���Q^��[�3��a��.�#@���R�G���􅔞�����<�:=�_o��ei`4Qp*c��"h�ǔ��\{<�Hdc-T�u3J���8��;�B^<�'u��ēy����u7�[𰬰���I~�Z���0�bo�xfi��3E.����jy0���I/���'b��-�ߤ�F����,�����!=3�T�9; ��~�ڇC����^.!ų�s���,�xR�!��yP����y�x����k����R)�pP�詰��R�˛˻!���\�Ouy��5%�{�L(�?��)uL<'�
��$�Չ���+��,��l�� gJ�*���\>,l<�]3�'�K��ӴwH��8��Q��15�/LO���A>��fӓ��B������vug��9��Ѭ�--8�0^�t�.[�1Ğ72*qg����x�bɥ����9�Z��gơx���Y(�G&HkV�c��i���蜧Y#<G�4��f)GfH���	Y�_)��������f.[v �ΐ��ĶmzQ'�y��&�Y�r�x�Wk���L���}H�Ϸ�8m^V��a���`�4��2���mskp��Ӭ����r7%dAET��F�5��P�
�hwx�򦞙r5�
&� �zC8���
�"m�O�`pF�\l@ �G8.ն����JB	5�-W��pi���e��k���Tk@T�PA�:��g���gT��	D��ϲ�9�4,��GV�`K��Zx?Ϡ�}3���yu�:T{�d5G���r���v
����0:y�����Z��3s��=��k�<?���WH���l�]�I�e��/T/����	�PQ�f��^ .�S��x�c�߃Ɍ@�X��bf҉skΛ�(l����	 @d��H|�-i��lX�S���Ȱ��������{L���w)�h��.ľ&���+?k���Is�K�������%������F�H��!���"�lDZ�_
5$���l�o�%°�/O��NX2����/���\iu�,�qC��h�\K��4{?෻�/��(�Mv{���A �����|��#������V8�����
��D� ��h���/�o�V��O�q1*D��(�|������zQ ��!\��%f��X�0#���a�iO���ΐ���$��]��#F�,)�J>~ݒ�ys�fX�?�iV^�Fy����+w�-���٢��K� D�,
�~Ð�VU��OfA��X��Bs�(��u��/WWt�G��M��h?;W��7$B�|�޽Lz`8`I���s�H�?5�� _��Z#Y���|2 ���'�662��q폵4���te�9���e.:h١M�Z��C��b���"�!�����lEK�+���[M�a���64��h�a�N�T�xϟ�Azw=*�w�;�C�W(�������L�Ufb������~������d14�N1yx'R{��� )a���^�dƁ4+�#$���1��$�����:��D���z���E�6���pqO�gs��v�_d���/4�as3.��G��j 
�6�r�~T�]�%�c�/���}<�_��*5�,+8�<+
��9�/h7YV�@"����<�co��ku�[}����1�&x�ߑ�o�Fߟ�j��`��V�^���ЋtQ-��� /Ys��:/��T}�M[�κ3.
G�N�*�E�@Q&u0��������������:�k�U�8��NAz��|��}`�lu0�Ļ/�5覯	[��TA��%�¯JY��JO!�(m<����9��t ��V+�1����ks�mf�vV�x��m�>��pK��o�z_T!-���U���d���<��{�oY��A�([��4�	�~oo���"��3�jكk-@Ϩ��G:@Ԃ�}樁cb*[�^�|(��з��|�̢Ng;|Jz�3_o��<|c
���Q�C=�b!��Ocd�����c;6�/��|����:$��jGjr<�m����ܖ��Vܷ1���j0aN�3�LLb�P���3[�)҄N:kZ��҅��Y*	H�O[5v���'�d�Jw�"|$֠��aC�YGr�_/�#��

�PZ��_8 񺲨:�;���zɅ�BN��A��,��nFn��9�\��d<�)�݀�v҆��*Y��J�}����FfA�Z�>:qyO�	nN��hC!�z������ch���W�fep�`1}�<�T���C�	���{�!��w\�$&@�iIwB��m]=�É~�p��;�r���(����Qo���e�[7{y���j�8}E6+ ��l���r����I�]2W-.rf��T6�~�Y�����G=�r|��o�l�$��;�-�s3�jO�����}@-�aaLVCಬ����&�8r�B��z��|Z��]݊c���Y
p��j�ң�6ր')�E��_�F���B0x=S�!���K �+�[����� b`I��r��٩	h�-��o�+�β�?z����3���0 bB!E��ǩ�uʅ�s	��z
��lҫʉXn��a��©�ޏ���Q�J��.E�@i�N�?\O���6�I#`5Y@�a�r�)�`Q��_�=�����Tᱎr?�W_��y��W�y'ղĚ`1|���]j
\T֑�i��������a=���}dC��u�N��#����//�2^]Z�B��g�O�=9��ْ	���3؁9���a �@Ӻ�`� ����_��43҄p�Ǿ����ƈ�� t�TG��7������VN��14�99N����ޕ���`(�Ѐ��F�-@���J
�5�q�O�M-�-|�K�4t�񷰉>"�D�W�%�(����X<ׄR��[�nƳ-F��Xr�Ы;B���S��G���+�#߄M�c7�Oaf�JbW�3O�ލ����kZ��b�q��:�05���������䅶-1n����,�e�z���hg�B�yy���H�IHMw�r�w�N\�������pf�Ddjm��U�&�" >�Ѐn�Z]�\�������:e��r 2�H.[wL�Z�O��k�%΄��اa��No��Q�����:�ږj�&QB'�;�45���P��O�ya$`]0V��㻉h�D�,F�,�0�n�I��ϸz��̠q�6(Q�ߑi��EOHx�%�Z���o��C�0e#��OD|�;(�(S2Q٨��W�8����m�XB��:B�ّ��8��E�ҟ�+g�9C����YJjl��H0���	sAc���/c7��x��i��h�7Q�K��y���%�vye�f��L��[�Ȳ�}��/(��z�|Gm�C��5R4�d�TޥH��,eׄYz�,�D�m�]��"Ԙ�&���0�c�1i���TJu�P���MΟ��o�"G5�yX��s��&ZJv��R勼� �)E"�,4=hY�g����!3A@� ��-��ڏ�z�l��"]X9w@Ջ=��dM��p��F�K��$�!�/ʀND��T0�)Է�&�&�b���R7;4���^�g�ɲޚڔ�X]���*��i`CX�r�#+�F�&�͡)u��dS��$��[D.6Z�%S]IL�� 4C�k=��m��䖒  9����t
rb�%�5���%]���X03���Q,>�z>q��:ʮ���U���7s\��#�0�T�z��x �*ސ影k��ī�):�>M������e����t�_��7e�Du�b�Y2ֳ����؜Ɖ�S<;7 �/Жu"�֯d�1��Q�G�R!a�1N9+w�7�)N�>!R�}#	\y��P���t�I{p��lm���q!���2�t�z\�S����r/æIC�d�Z��/�����4�cZF��m��n`�-b�E�^�]����4⸷MF T�����)p��~�mV��ժ٤�o����Q�K���[d��y�S���Ư�h�41 x\]5� ��ys�N�������`�Bc�<�CV�\�p��p�1�3�o%��u�OP},/Pf��mi�Z��U�5�����tUh�!�����ng6�x��1C�ZCMO ��4
�&[�ߧ���F��B?`f�BPW`�l�J�e�f�9�6Y�i7�.��&���I���C���)��m�hҤ��ܘnަ�Tc8�*�R?���M8�������/I@�sv�c�+Ay�BB��ђ���S3t�b��<V�❐�D۰�'8�qL=�~�~ߠ���Ub�C����c���/X��8��8�M��ĹY�KY��G(�'dH�7��u���>��ֈ�?�G�� �A�p�z��L|��E�y�o�\*��"���6%Su��O�4�Cf�H�m˚r8J�;Q4[��W:�ܨ�4��5�3Pr��������,4�wxX�g��y9"MGHi����0��En٘�(f{<}�ݜ�tG����(��⦿6:�U�/M�`��}��8�ϑĴP �K!��~_+w���v�Y9{�/�J�a%�� 
���~�����oL� �+�n�BRG���@=���{����F�;$Y�X��������4�`R�������sȝg-��N��u&�

l���39�ڢݴWe!"P.[��N�}��^���o�5�e5���a�)�;o�S��'Um�ߗ+�z+(�E��,U*T�潺/�ܣ[Qy���/�
��2ul��@��@\lW(���KQPb�	E	{�RQ2[�i趋�ν�ĩ���k;G�x(1;���E��؇ЈE*�1�
�
���k<�$���+C7:r��J/��2��7��䙩��k�}���>2)��̑��.d��&�I2E�ڹ��%B��q&��J�}>̰����ʜ�*�v���c|GՈa�S�����/��H��~zZ�n6��T/�/�V�`��B�Ŵ&��j#��0q�W���d8ƔJ��@� �|�%�5���ۇɵ�Hg��	���h9{_��T�4GLV9�f&���A�F����5�*��RQ��3W{�9��+?'�(!��fུ�4��w�=N�