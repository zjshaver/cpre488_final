XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������Q��z_w�Lw�,P��!>���]`�(n��a��c\�]����P�?b��G�$�&`��pQ�8���!MԿTX������l���js>/0N��ZDg�6�LM���a�L��{�W�8���X��5���9Y<�N�����/?�Vn���5l�7�Hr�d8
d}5�=�"�z]�ꬼR�ﭹ���YgW��Q��7J���sM~��4��Y�0%d�wo2*��X�V���OG%�м{F_�0�Cݵ���x�F"�����\��-�p{hi���	0�o�g #���/=�c��r�|�:-� �Eﺐ!�>Yh�Sqq�C�>�����a���Q��cF�[)}^��zoe
U�Pry��M�@,G�:,��5έG��N�n1��C�Xң���{��̋�jZ�(U�ϧ3c&QLIc���@�=�jˇ��y`��J)����Y)=������(�"���a͉�Zu�������椰��P�'eq�_\�Iގ�"?`��>�¸� ��]I9�1���c�|]��^��Z�p��qSK������*NM�����~5��\�9�\�Se���$����L&��A~v"��j�1N��8YV���sq�N��QW�)�%�'+�?���:��7�Ae���<Ę�u��
�w���Ag�+t=\�W��V��c�:�sX���o��`�b�Akŏ~�8���.O�)�:�\�X�`J���	�vv��>����Zз�Aߦp?<d�u�4��XlxVHYEB    5cad     f00��
����%O������| p�'���թ��\/�-��<�4�(q���%�@�l�$T�kzd�t}����#�o�QP�f%d��a�I�T�#���|��hO5�Kچ5z��z���2.p� :TT�q4�
 VE'ѕ��U�[>��4U�g�tǴ��T��'
�a+r�-����)��|:�~%����K�`\�]SӶO*"�N0�ߕO
\l՗���~����̑3��'4���k�
�3m7/(���x%R�2��$	h,����vm����J�p�0������\��� ;�$�lͲTW�lq�d��s�a��qC$γ�cw����_�1A�����x�6`��*�agJY�:��uHyQ+�\�\M-@^E��؆O��i�����IH�o��Ju���lN:7��W���kgL��ki�(�٠l�B�����Xn�S'��!k$�A��R���-Q��Ok\,����×:��7�'��}�+����I����o󨍖��S�A[������4B��F�^��5����ߘ��y8�L.�WE(P� ��*ҏw$Y;���%�':�-�t��W��w,��ӈ�ܗ����D<�@*�w��<��A�n�MK#��*X�ES˰c���B79�8ePP��ų�d�J#}�Ű�Oz��m<�L����pu�Z�oǥ� J��w��k����ov]�����mޥo@'{6A�����q,�7 (��h�d��wÿ.(�F \�;�y; �@	��;&�RE8a�����4em
E�50�`Y��r;W;qI��6t9��0����`لw"���Q��Tl/�>摀��s�I��lS?��ǯ �Io#]���l��)���$^�gEZ����&(<=�FT����mG�Q�.j��B�e�\�H���A���y'6���ìܝܼ=��=��14���v��Ŧ�(��K�ɝ�x@>2u��pQE�3Nk���eo	{�,��֊�\w�T~*Ӝ� �l�0�inN�?R�QR׻`B�]���S�<q���gi���U,�`�N����BV�`��J$[��&������U0�N?�h,�͐y ���=��J�"���oWC�]l	��߽|�ۯu2�zD���^�8�����b�9��}�%�&�`�Z��t�r)*.,h���_���Y1���*�D�;,g�tW�� �	�qHO$��}� ̷	{�0�>��r��|�Ǧ�A,�'Ľ+_I����1���_��2Jn{9���y��+�FP�L�~�U_"���6�͹�o2M�o_��{ �z�9�]���m���&�Mo�{���ޥZ��BūZ&����ڝ�#D��&o�N��k�7`��&%]]É��^�7��w�I0��6w';c�O7鳌���5EL�������^��Y�"�l����*����$���N��F�ϟQ��y��"�6���"��tF��
�0aDe(_�9�x���g+N�����A;X��\�9�� ������C��W2�#j��*��r�E��6���@s%�FXk^���ȱx�2��]H�R�P�+,0YI�M�B,>Dx���TǴti�}��|y�\�V ���W�!~��w(�y���J#�É�܂Ge�.9p�DY���R,�۳9�(�;O��E{�É�f>jm�;6c����Q�5�-O/!Zbݗ���_��
 ����l���3�'#�h�S�>�{�#9��&Ӟ�׵O�c6��N���Ź/;�V��I�y'3é��I���a�@g�"��A��"�5|,.�sjr^܆����qz�����(i;����x:��k~�ga�p?"⼹���y�^ct(�#�a�K]e��Ū�Wt c�����ߣ����P����0���J�\rmb�6���s��?Qw9b�Rs�^��捉��Hs�E��t�c�?�OAѓ����c���ߦ1B������d��i&�y��?�f�\�P���B��ٷ�xד������T���wǖ(�Z6֥��۫殀<��QNL3x��s�ț,bJ�r�Xi���J���B�asR��x������?���	V��?~�����w�Z#sv.�����-��Da��A2�E��oGl��0��Un���18_�\����N�3WlT7�?�ZM6Wj�:� JuP�*��a��~�sh��Vt;�J6H�<Е��@���s*��a_�B���rb�
��D�&x�j}E�@Q�Cn��hn�jGC�,|=V�#>Up���Χ��T;��3k�i������Ɯ����?��ͦ�
�Ip��&1���n���K��m�(��Ǜ��c�0�(��p������^�m��	2�͍ݢ)�i�#q�W���Άߊ�����Ҫ�z�cl����pq]�ٲᡓ�hչ��j3RIД��	F�Q�N���&��~����ߌv�4�}#X8��=��E !y�X�s|i�����?Z�r�}�h��i��$eë$�Y[f^W�b�^�Q�/%G�]�0 �.7[Z@��L����q���gm�C��%��o��Cx��C}:K	_2�}`�\�6�Xx)M��n��Ή}�A$×�2r�c�>�Q��Y5�h���U`�.8�5�>[ŮwˌyX�
��"&�l��ZA�n�䓬T���%���u_��7����3�|��;�g���D����T�7�t��.��jW�!�&0Y�TXX��y��8�����x�7i�]
�0A�٣��Ӛ�.������j���td)����q_ E�̡��U\/t�	wJ�=Kg{��TGH'pv���I�ͣ}Q^@�3H=b�E;���������J~W���G�T����a$O�*UbCS�G��M��oۗ�R�W,�J?	�1z�Q)Y��LL%���1���>�E������oמ�?�N��ٮ7��H/i���]���^�w�SK8��t�=�j1c�/��xk��y�K ���W�l�@�i{&ni˞ج��b���&���T�ǳVx~l13�8�I_�?āՂ|��w���`frp�� ��#��/�;�1�~у�2�5t�!_E?�z��s��¾�N�*u����$������U���v|pa�>�{ŃɵݑVCb�yu��� ���U�8�vO��&gE�����,K��R�d�}��uŽ���Ө�a�`=�ey�\�<�7Q�~w�-��8�"�RISIV/��U���}-hJk�8����#ڗҖK��X���
K��C{o��-���{jk��J�%���J�yO�w�t_��R����퐡�Z�p����p}$��K�$G#�%�����۟�#����("�m�4p5�0o�?��BT�G��P�ܮ��
S�}#̫�����G~��/�H���)`�B��^���}����iɋSp�F�x���HI�o6	7��w"�B g��uY�Z�e�ӰT֒��oCb4ߝh3��\����Pw7�;"��A�B��8v��������%G
��_���'#�'_|��I�Nc��5��E��J��,��Bհ_�\�g'W�빙)|�Ř��)�Ɠ��:FG��LZW��3�����p��ҍI�Uȝ��]�1���&q�i��HZ����i��h؄�X��+�e<��x
^���������מ���J8����<O��K��!�&`�K��H>Ķ2��[:z�K��bZh�����m����Le4��3��rqL����� �<����T���H�:6�F�?�\�|���, �Y