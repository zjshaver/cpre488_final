XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����tL�2j�$ խ��f�(l���4�,�� �ǋ��q\�p�V�:���J��2��b�J��ӳ��W�W8�`\B8H������y�4����gR����{TCD�顓5�����R)�7�^��Cq�-
~|����i2[�	T�lT���<k�E�rD���96�%�Qf���˲+["I5��r�qX�9������PF.}�Q��w]|�e�7e'3Ng�#��\@��G�R��4��ˇz�0�����qN����	�S-�?7�g�L1&�����_�4�Z��ΰ�XG�yƪ��c�K85	㵒���>�/|Hr���Ba�%���w+9Q<��TU��bk���C?h���!�W.��1'���z߀({�Cj�Vڄ�1�A�6�T��p�G�Hڳ��8�:d��z޿%XW��"W�2s��9���&�|��٬lZ2��%i=��l���.��xE��C���$K�ˉ��
�Q~F�NnG�2�ӄ�u$��k>>yP���ӈ�[��x aV��F�9�����'�A-_ܮ����<)%�=PkY_�&Ԍ=�<��P�*������٢��������GLg������8�[||�R��Z>�8�Tg�Z�%�\�Ϫ�e�zh���y�$ز���+�n�$�ty�'8�/߻��6	�!�求.GS��n��p��-Cpя��Ϡw61���z7�����h`��� i�&�X@Ҧt���LY*�fS��Դt���+��a�5XlxVHYEB    3d43    1030�^)�x�Y�o��j)�����cR7��+�Vﲈ�2��V�E���u�=�k��N{Q��W$���0�1�/l�=�h�/�{�e�iO�o�k޿���k��,^5_�_3L=Zt�w�m/���[[]п�A��1M�� �q�c����ˢB��� �Z¯K�R���f��N�Cŉ=0�5
�a�F��,7rK���箣zcT$���ʫ3�sO0M3Q�O��Y3��^EV�����[�'�g�4����]j�	��u��H��s��*t;��3uq�	?G�S�����xc��2�a���r�f�������]���̎��#�\�ٗQĹ��d��h����Br�a�*q�?Sl��N�q>#��?���W��� �5\�a~p?T<B�X�����Fmt���O���� ��j'շ���>@��P)��[$p+!��}��C����,�j��׵��v���wJmHX����I����}�*�8j����@EQk7c�'�#S�sW�Q�n����ȐXH��O:�h�W��4C6��/�B�9TOYL��bW�����:�7�5:7�������Ӽ�����pߧP�	}LcuW���䱃��<�$Z��)ֶ܀
ˮz!n���/���U˱T]�cB���$D���m�y�}�Q�! T���Hi�C�';Ҟ�h�n;����Q�Ŗ����τ�G�h����t���H��|L̈A�
�Y�	�{=Z����!�3D罵W�����K t�_�a�{�d�B��"n��K廕l=�sT�~?�V�0������vQ?���z�]uGh0�<�����Rb�[\x:r�b	4�-v�͆0F�h��w�R��r�DM���3����,����=�$3�}�o��{��
��A	u��vBE$4��1��Ѕ.(C��f4���u~�#i����+���JM����r�Q\N����c�u�.Ф{ͼ]zPU��g�O�~��IV"q��J��d
_lR��-u�/�-~5@	'q�u���Yk�(�BV#�9R��{��kaޙ�qveSiy�ݛ�O���g9�r	���Pu�������+�~'Ƈ󍕰Ƣ�Hb��r�%��j�"������W>w��$6���Sh�օ.@���ad�p}F����M�=�n3�d�d��в�_h\21N�8wdiʆl� #�{Ӄ��4߰�c���k��"����NȬB�F�צZ�S�m�N"��X0W�ׯ�2�v�Z�N�#:*�yE�T2H�J�WӺ��ˬ̬��x�`j�E�ѱB��ٴ�0��W<���^�vg���ҭ!�E����"^� m=���|(r@v6PBޮ�e|��=6�T��)av'>xV�@�ւ��>��1/�}D����͋`�����\�</1Ɛ{�v鲨xp����Z+�5PPCeP?R��8�|���,VV�F2�x�Ax�ZWg��x[���g%:�& ��/z��w�{�����9X��3g2R�X�h���d����(�-�I��%ە�NE��i�o�țj���@.�h7���&��pQ�"I�L�c���lM-�H��xwcG�/ �v��A��)J�,u:Vd�v,�!A�A�c[��?�a>ɹ��S׋|��e˝˒\�k�S�]ͫ�_W&�J�Z�bc��G��5Q���ϲm��0+���N����M��U�y�F�r0��=um�nVk�5���X'��ٙe=<����ϤY1�6��X���E���]�K/� �ă��k�ꞹ��K,qn����z��{>�����!�d�}�%@L_��t���nͿ��@�"���Z��=��S�1YbUk�Lԇ=�):qD��EH�#sח����Ĉ�0���rF�
)�B����|n�Mw<��@? [F��a-Hf��c�;LTvk@;�։����Ș��T���� �ag�@�)�@�����#z�lYe���;�|�H��>���ݛ�W��X
0:'K��v�'tʳ�#_�RZˬ�t(��Q�o�R�%9���[�w�i�ܖk�N�4}���S��2�n��x/5�<��T#;�t��~��8�o�r�ڻ�Q3*(sx�?����_�={ ��ppbu�E���"HtZ1Z��\3���P�mD���U���J� a�%&��
�_5@5�F�BFJsmG�uv�[
ē��E��ƅ~��PzX\���i��\o���d�b�t�)��~�
�_8ǐ=R9g��Cbex�^� ���[n�ۛ��TH�|]jC+Gĕ��Ҕ{�G{�TA�n�#�$�i��d�lѬ(�����$�>.	��J�~�s����-�\��:��nGX�A=�,� �s��d"��Ò�Y>�l��_�0 ~� �^�3��򥷞�#ܛ��@�y*�R8�/? �B�e�a7��[6�>��z%$�Y�4�f=*[��)v�Qx�pW�&�G$�q�N���\���[�!�ե[X�R�2�{��uee;�ۿ2�d������J�Pp,�X�@
��jZ$���={�+���?2�64B�Cs=���=����M󅖬�d2R��ضA���룵5-/B��U���� �C�n/~.XX�f�Z6j��~'�������B!��7R�-��JL�S^�3Ӵ�
�H�;���]�.�wj�
-�o�F�V���]�B��T�k��~P,y��$T�ߍ>�N��̂�.ڐ>$��Ի�48������f��V>��R ���)h9�6Š��X���:74V�ȕB�e%���cQ��^�����a�~C�2)o��Px�
��x��>�pnJ��ˋ��ΥJ���=�1W����&�x�a��fP�h��������	ZC���Y��{��$XE�^ج�-��yK%�h,?{�5͂���L��j�I��^R�Ag��=M�h����,�!G���יpdD@��U��|��@��z����&1N��V�s�H��Y��E,&˗�#C���;xH����ɳKd�{N�֏jp����%o��� C���P���,�,����l�'�wĴa������^�E~�&M�=���[���c[�V/D�5�׵��\Պ�7&6]ik�3�e��ϟq-M��۠��2��6Λ�0b�w��8N�r�dDw��:�̐Q�h��4�Қ+�HS�ޡu3e�
/�D���)���@���寅}��v��f=F����ձ���Nv~�`��+n�ŋW�����i���J6��ج����T,����� :4.��B	4��7V�q!Ħv�pe����/����X;�R=���p�D���հc3n��U	�v�+W����ƽu��7Ne�U\r�9i_3N˃���ɖ���u��y�g��WUw2uX��vz2��6� >�(�Qu�uAs����Q{���d������n,}��� Ϡ�d�
���]�}�Q9<|\]5���s�5�[A�ʓd ]K�ElA'�Ö�ԫ�j�1*�v�v맄Y�'_<�z{"�6�g��ew@���p ��ji���;�	�֊ ��4�3.���*=�W���җLX���\tw�.�k$�bx�ue�)�@����ϋPzF���"j��H�_+J����Ί���vY��ă�ReN�U�m�2N�L'�%��N|� "[c*�Gbg琈8(�6t��͋���֍� �͠��[��N�١+[�-7���Y����Aq��;\�w�R��Q��x��z��M���F��u�����%�w*J	EQ�)X{�SLOѪ~\��Yk!
y��:�)<0i��Z��o�G�;V�8��g��bp�\�M�2Ԓ7�$���T�I��tl��Ő���� �D�f�]4�� [�jS���5��#�q�y��=1�ޮ�����\�����Z%��J6Ƞ1-"�㠭Igp"jL��/���i�C�^	�'^�J2ci^����h�I��`Bc�!���[N�\,�E��-2�c�e��/ޕ�ɔ�}�t�5q8���y2��"��B�v�w�c�2/�QN|�5n{+9)������g���d�gI������	�\�r?�>욎��X|ĝ���oF�ý��w#9���-��C���Aˢ4:��.0DGá���ƘF4