XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����ʩ���rM��)���D�jG�?�	�{ؔF6��~28^ :�L���L��;���#�V�<!9�K2���?��(�F�!AH��ЙǸ�y@X/����a�u�;D:���0��_k�������d�	��-���J#$�]�U�Ɇt�4��vI�<gP�֢��ld�E�D���| �RsŢ��T�aK��\���z ,� ���������?�`a��T��N�mI۫��7[�Qx��X��x)H	Jj	���9{ROXtQ�9oU4��� ���r�����\3�^h�V�������j\�1���h�m�l��$jK�8�H~7��7b�uMABݤ����w!Ϩ��e���SEP+�B�.�:EL�ְ��_'!&�h�y2��S��`&��9fr��j �4� ��i�W�Ӡr,`��2���lJӼ
wP:�&�  �w��#&\f�m�1��F[��	p�:�RI�i�G/�1w3-/p���\� �]�R3�p��KKf������D���=>�g��Y�B���8��'�u�2�)�r����Sd;2�(�WN��l5��Vb�����+�v������k��w�J��a�����t�Ȱ���֍��Rza_,�}d�e|c�њ�Jse#[Z�gV���G��ݵ�}�M�Z�(᥷�.�u$�w ����Վy����!A�縥\��8[҅���D�����?z��ſ)�p�[�]�J ��4d8��x�;G|�q'7ᤤ&ޫ˨*�7�a���XlxVHYEB    4052    10f0��J�a���Y�YM�g
_��O�5����V� �u�3���淪\h��6��c��,BLi����eB"0�!�RG쀇��n����iP�%����?^��V��X�C������}�G��_�����
��e�״C���j 0+�spP�ξ��yҶ�	H��Bn%��\"sp`�()�ԫ5L��B�L��َ{R6�(@�m���ݘ>y�Ni5��8M� � 2���zCx�/o!O������"s�E���^l�Mi�ڀ;����Q���Y�bF;��N�����dNa��g!s�>�z7�[xCZ5F�뉿��~�c��$����"r%����Be®���ܼ�՚II�[�*�=��L�-ϧ ��ج���;�Clbr�]��Oa�<h�s���ǻA����a
2n�J=�;<��*@Ӹ0P�!-�ldsU�/nSc��:��S�k���.H��؀���v	�C�F�#�	�a�X��D��#�#��Pט~t�0��'PT,�yz�dv��u���"V�Ϝ1���=��D�|�4��i�V��{ե-*p���˘�1��Oq��u���T�{��a�4R�y�d$D�����U�8�wʠ�.-AX�@�;˪\$�̶>B�W�P4���{z��R�2��?�ZޏE���I�	�II���{R�H�dG�����|"ᵩi�M��d���2�o������
g�J��[�C4��:��6!��%	����T�x�� �\��O_F�Qj���@�E��)�m��~CZ\4]�*Y=/ ��^��t�Up�lv�бY�1[�����Ω���������5iM$���m_�����x�N#�}��k��V�F5�U�M���)�a�ş���$��:|.76Fu�#��ˢ?�8��ŝ��Ϡs������A�Ё�l�o���H=������>�i9Zbd�Е�"�y z
z�U��)�0f�9����k�c��6U����7!��n M�(x`�� �_Eb]��}���u�Q�,/�����_߶��M�<�΅u!� ~E�>8�_!퓵CE!�i��8��jhQ�o+�/u�e11Qe/��0�������-�����u�\]$h�X�o��_Uʍ�'��J�tS�v�`u�V۟1l��Z�rBFc�u�T��}�9�E�G�ߊ�'_�P�3eZ<�����*5�;I���k$�w��ok,��Uw@f��_]�b���@��n5��v�C��uuM��5�_ouˋ Q�V�>.%m��!�$thHz�
s>ܥZ� x4I��r멳ه0��yl���%b�)x~4a�iО�@����8)uTV�m� �fc�o]b����Sց'�)��__��n����G3c���4���}A:=�+�r�� �M����֨�#�L��8J���wHWW0�g���<�dVL�������;N7�nYpmnl1}���m�H�yB=(�D���ޔ`���f�ӓ��GLSs�o�� �(sR�k��z �O��/T��i�j��A��G�ǭ��J�X�p�~帩�����L�S̺R����+׭����8�U�}�U�H��nT����5vL�i\bK�Q�Y}Ks?�����N�K�^���0�Ay5�(��wf��&�Jt���p[���!w�u�L��Z���V���,�0 
������Q��N HO�����*�^D���^�&�) �i�Q������-RRo����No��.Tv�q<�c���Đ`�-uQ�>�E�H�j?0�0���Zo�꯾�Ə�n� ��H�>�^c�/!=c.b�:�T���om��87I�ٴ\��N!0C]�ϟt폾]T�S	�WJ�#��8�0Bsv���f]�J�|��������,('Ze0�'�6/6��	�m~��@
�g����VM�w^�ޢ�y�<P�0�+���G�c���ho?��B1w1�/�4�yq\�r�m��3�<��U�,��GFZ��r��[���ue��4�7��+Qàk�鱱V����l�ǥ{���i/hg߽��o�K��-v��B�E��v �x�#s��9�>���I&k;�}�v_��YS7sU[aرІX�:Vʐ���?���T�qr���l>3@��M^ɟ��0�d�G�����Ӭ�����GZB�.���~+_����YA�xw���������Ȑ9�2�xY[s+�i�ϩ/R��.]�.v�Rᣌ�*@��
R��6���V�F��'C�Br��R��ŉ�e^]y��s|��R)LDg�_MV��-�|BV�j
�m��U��N��Mv{͚( >����Ӌc��^�7"))�/�U�k,�>j�U���2��_�_Gm��
�+]-*v$bz�A�'hܦxHG,��	��e�->�B���P���[w@��f��,����%3Ҋ�V3<�#c�E��R��tm�j�9?\�vk��ԃV���h|3�h�w�s70���1�0��	y�o���Q���}�+��/��,�������b8)Q?�^/��z��Nf茛AUS�j�$$���SI+��&<��J��˿DqoK�mPǌ��NGuy���� ��L�/(�[1�Fu�a���׾ݳ|A>�߮�[>�b#ތ8��AfݾHkL��%$�+(��5l�'p�\�>��Ei�2h� k���.F�o��0޵ԯ�R�ܻ��{�#Ft�m6�¶�LĒm ��+n�I8���;ظ�*�����'�z�$���e�����j�ű&�}DCe~�XQ��I�R[������xպ=度��]Ǝs�,y?�b��N���Y�VY՝i�H`&�@�KqN�HJ)��Iݪ��-���٨ߊ0mħ�����)_��ٟ��網*�R-��D��iI�T:��h�����
SP΄����"�:�ݨx��wK;�L����W��-1w�8*�T���������!�ٗ�l����U6i�:�T�${�:�	�$��$����'=�F͠U���]�k���$;�^dq&ӝ�����K�LW���a�J�5� �e�`'�HF4�6~�m�ͅ�}d���[5��}���MU�^�d���>�O2O���銽-��C1lK�
��1�tM�`�S���(���2{�e�e�y�a{[� Ρ�	�����p%_��hߗI;s���ͫ}@��!�T���6zB��IC�-���f�X�bsE�I��Ldho#���%�:�k�l8���,FoJN���\^��j֔���`�Ԉ��Z��NV�Ɨ��8�pC,hj�F�h��4��`�z�#[6��/B3��<rQ��c���,b`�A��f�9cLћ�TY�{��W���1���W����ˢ���dƔ. �}J��w>K4�m�U�����?Ny�,B參�

cr`�� �g&1<5��~��D�(,�pA���wܛ���<��ek�b��f#C�>�hk�aT>N)ǥ�����juX�A�� <�O���~�:&ܕ�'���kj!*v'�!�6�����4�&ے� �ޝ�\��^v�a��9�,�����Aq-�v8�e.�^��.y��7J>�J���x3U9��+�)�y�iA���S?��	��1-�TN�ʷ��X��5G�c#Q''7&��:[�{3���Z1�j �y7@���E|�ܝV9�HC�}LCNp����.��R���w@�
�{�}�c�6T��N���ʼ��Mz��P]�P����)B~�]��qT!?������c2��*�@3��<��o�0&��8����Vw� #q���Q����O�)vec�h�	����� SF�>/�,�=�ZX�LM�so��ֳ��9X��FE���%5ނ��^��x9c�R�O��Y��j��=,�� ��������Le�1�N*�S&:w$��Q��U;���ow���@{ֲ����8w ��ރ���������v����M.���o�C%/nr�U���23c8��R�?Ʀ���+�.�9����;�#��=���6�kפ���e�p�	8�c��.�K��R\���~>ǣ�eA��>�	�����g��M��D����#ё��f^�8i�~�ϧ�bB�|q�D��x#������R&�Ĳ[��5
�WgzN`H�9��r�.�R|KN/�����q�M�w�+�U��*ɨ��A�Z#��@.�c���ҡW�U�7%͗@�v��&`;u� O�w������[Y-�������h���>O�%�����/�{���&~|����]�.��ib��p�ߥ �J���v��a��l��z������	��/wp�y�oi0@f@3��I�cU�e��f+"