XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��^��a��y�]	�A3�;�¢��<G���'���>&���egI8`�h�Y�)�� ;GKV�`LE^k>���u��*ݺ�g���G��?eN��$Na�w����߆s�Xr�_Ldp�So�e�UN$i��X��N����}�`5Z����fA���G�V����a�u�}2{��:tN�8<���j�xr�Rʳ���U{y�)o(�� Imy:E��:7�Ŏ5�dM�n�f��A@���%��SC����1�@�=��?@����d�^��7����!	@�J��%��N:H���|��h<P41_���s��7������h@NG���m6�y�6	�K���Q ��0��ŝɹ�Q�	��J�>���UU��r�$���u��s�V�ה��fNy�ʂ}Hy#�B�PؑM�i/�D��#!j�H��H=U1@�3ʛ�Ҿ#@�=�mB�>Vٍ�����En9�Jj���|E^.� �#�Vi��4{�O�th�4�'as�;��e=���#�b�j݁9JOB9�T,G��z��P���R�On2�X�v�v��^X0�^E&ߊ�2�+��77 ���[�T�8�utj�=��I/U��߂����H�N���H���E�ӧ+�J����#�誓U���t2����Ah�{6��Ч��]ꚭ�;��_���z��+�)�S�����V�%����������}�T�)��T�ݽ����;�=?t�7'
O��Nw���v� 
��nm�~ɖXlxVHYEB    1847     900��	����w�H<+N�x�@����*���'N���p�����D[�ih����0c��K�HH�ִt�L7����~CxΜ�Bo���8���`2�ٝ��!�]
[�h�kO'�
ʉ��خ���_�<L��U�LW��<��(��8f�ls���)>�I� x�|�_�֡����c�#(��7=B� R�ԗ�@�҂��f:� y��g {{�}�wz�:4'�['�p�mQK���	B�]r���7��A�ElƳT���i�\��ml�{lw� [�`8@9Ȍntݪ�k�ؒ���5D����~�
�*��"r�/�7�+i�f�Q�Bz���
+���\(Eph#��%�>PV�?
������oLK��Ƥ���|�I���`�YJ'���u^򨻲����L����I��x���
m��X���3���J,�%�A�s�	�<2���e�R�iQ��+���!��M<�Me��%�W��\i�6���ȼO�����=�!��6!H�Mݙ׭e36��D�-���%���t�2�|�B���� �؉����C����|^�2����Rs@�7�Kau�l�����ySk��0�(���g��aMOM��J�	fZ�a���Ȣ �W���$��$͉��L1Nl�;#)��N$�j�e��kѭ���x���� ����#Ȟ^�b$#2͘�e��,',>�T��5�EY(9�V?�����'W ����g��A���u�W�5�{�'�C���r��ᶵ�#��6�
�;�[&�0�X֖�4�X����<�u�I���NB8V� � B�a��>%Zj
t�¤2S����A8��5ǯi5NU�8�&��8�	*mb)�;H*�pm= A�ɵ������g��XS/}ŗ�����J|}wVu��z�;�V���O�X� /T�,�S_D��2���I��N�3�m�,65&�UBL\%qSR-tg�G���c�uM.3y��a�����=/.�Q<��Њ�~ֽN���$�C�
*���w� Մ��<�	����:�i|���g���f�����8���a��v!"Ko- 9)8
�g�3Z�OD�����ԶG�O����k.s='�y�f�V �)�fɃڰc��������'&���u?���	��z\P�f����)Z���0�<�{o�G���OJ��Ǿ�wfpj13h�XX�WA+��v�350"KF���N�u	������D�^]>���Fb����2�L+�f�N���\`i�w-r�_Xn.��k7�҇�M�k���S|^'����#=�K�}N��
O����С�)�m�mchg���.˹&�i��+4�Fw�+>��l<"m��l^�S��/��/n���lp��k�� G�/����ŷ�vϼ� ���#��ҧq7�����x3=,?���VT��h�D{�v^��5�
{_����J����uP(�732�"�#��{�x	���2��m���װ(��4jʲ+�frc��{������y����CKc��f�L8��q`?��4H#ՌƯ�����:/��lC7��&��R������| 
��8,;�?�n�f�^��@�h�!ƃ��*����D��Q߆����e�������i�{�����ƚ���#�[!�>�:nbZ��(:i�VTc�p��*���Am�r��9^�e GB���Ĥ�`.������	���DG�D�e���R��:y��*�y|v����X6H;{��Ud��g����;�=P�#R{cH�|D��Qo�_�P�x8 ��)��B��L�-x�
d�� �N��Y�9. �,�}=)7(q?���.z�}���&Ծ��o؄������T{*xH�
�x3��Gi�V�ټ]W��й�����6�� �Tӹ͌,׉���4E�Ꚕ�9wWJ�o95����-)>���k�!��G��T
C�)�-qU!{u0��g���n�T��X Am���Z��!�}PzV�aӢ#�� _q�Z{��!�Rۧ�k'sylu9-��J<�s��a�-S{ΨL�s����1OY		5�dYC�g�Ɉ�2SL`0X��hU0F���P��=�9g3��;��"��h���h@Z~���O��
@
颹��.cG��oN4�5���'�j,w�)'1�g$E-��릂	fP/ץ�X�כ��׵TYÀ~�I~Zo��vr�x�X��2��%��b��ipk^L!���He%��]jCs�O�!�D^xկ�x�Iv�i���C���i3��]}�