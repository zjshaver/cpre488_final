XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��gȠmӊN<�5!q��ߺʣ��x���g;���x
֌K��趗wv���
�R�2!��й��TrJUY��5"��%0\��1œ�s�r������EOč���J��!X�S�7P��Գq�V�V}%f������$k��K�v��X
D�1��O`<�+�����6����*_�E8U���������P��H�~sM�:/�*����gFhwb�Η����2�`��t�[؍RA�v	�\[ jP�v6�x���g>�R�Mq4���d���rl�S�蔀���O��aq.;�����|�`������_0;LfG���嫿�/�`�x�����g�{Cz2�IW9nL'���A,,?���9�A�K�����N�cB֗�)���v/L�HH�k�hJ�-!+�|Ѳ#�D�%��������_f�������Pf�阽�D"}�,X6q��>�֟�g�Oh6iX�C�Zy�(w��
�~�-�^��Hז� ʗCG�ʣ0P�"%׏;�m>������6n�>-*B��z��U��A�X3�A����jȮ�3H!�K��%��7�֚��ڼ���rg3�PS�O�J��g��ܠ�M��Ϯ5�tl�=���\�ܛ�9?�\�Bx3����D����	���d�*��=�L��
'wD��+���y.�ύ��s��,P<,�uv�؊�X��2�7p�$�����c=��V�'���h@56�_����J��t&555N��ξ'ט�a��hDV1}JXlxVHYEB    1847     900' �1"R�<|u���l�[�w¬ � Bx2ـ�U�?�q�:�o�K�x���c(�a�k������i˶��^�7f8{�!�Փ���6��sF/%�Ԓ��"�g�!�Vʽ5���y�ҁ�|��>V[Z+��{W�2��L�5����ƾKS��^�7U�!<�=��4!��Y�p����1!�A�H
� ����;�6F{#�]p���4o�D--�KԴ�� G�WƵMVܨ�X�S폪(�EI��i�3Ӈ���;��=�.�����f���<�{Ey�M>�<��uݱރ���^�N*a�#�	N���K�*�rӖ� ����z7R�A�83����������]�[Җ��L��2��p��H����[�b,#2�-�����t��*�t���%�eh3 ��M�����«���4�N�RS�غj]9�.�&ܛcn��l��W3ɑj�+�B�t.f7��9��f&,�����`eL6	`+rP��;��[�ú�Gt=��Fa�����Q�^�Zz�0#sX`/�' � �w_�~]��K��y_a(*�!��.?�6�=!�`�jgѠeI�OG�7]����g�e��C�ﵢ��������fe�:`�(Um*�Q,�+=�x��s�q#�z?�9Ű�D�M ��u�%��� �«�I5d�� 4���3#�q��g���U;�3R��z�/�,�����X��7�+k�n�J@�J4e��<g%�߷�`�K����ͥ���j����<�9[�Rd�����efG�e�c��>Qڪ�;��SM��yox6j����1�P���9�0ۢq����ye����	�W�	-��lg&�%��A�0gF��_��S�JȏH�+���dIP6GUP �D^���)���c�<�^�N�������?U:����0G
4ӈ�Hnf����Z��;N���}Do�'!W�ڞ:�9Wcs�Ҿ`��L�N�f�yaG��N���-'˪V9k�����wN��Ց�!����}��!ח!~rr����+I�j>N��۝��h�g��h�e����+�Q�ޯ�$�Ef5�1As���*���񕡯rv��>�F��eP�!��HHT����8�i���>�o3����K�]�K���E�����#�j�"�6�8���<`#�=�{���:9C��ӱ wG�C�u��OC�	k"J�'�ph ��E��z���T��,�7%nrjOo�qf�H�)���.��	\~���
���P(f0=}I8/��pq?�H(9	Ǭ��sم�F<LY�L�R�렑��E��b�@�9���B�f;	i����І<���z���<�ׄh2,� �M6�>l��8��bgvn(�7&u���D��.Og�˾�8�id�G��q1x&�a�%����RGfL��b��y,
�.*���&4͐�#%4�=*J���8��ޜ�3��S��ǔ�e?,�0	Ӯ�]p��ق-�/���n�?�e2��<�&W�SU�M�K4|����W��S*�A[yj蛣
�t<ڳ��)�"��:�D7��ӱ����p?�8����kN*[��u�zR�ի�p���J�H�a����14z�ժ��T���R8��q�W���d��݊q��j{_��n�8q�]� �#�2?��q^��:�5T`���E�/&�h�m�֯�p�H�I[����:��;�����L��eR�������ӎ�Co�<
L	l�!S=)B,�~��f��H�~���}�^�����:ջX��jXi{1pg]���M�+u�,�	����4+��i
7*M��XvlC�qv��4�����$Y@�эKt�0�J>�A�4ѭ�'� e�i��`uF5�5L�zi������C�4�Ú'JG@��0�A	��� @��i�� 6y��;�n��y3B��0[�#kN������z4�^��u�q��� 0��Z`�����eD�_�
�bP�����c��@!X$�^���U|��d����t��I��)���Җ�dH�	-KS��\�Nw��=cLđ����)#\�ܨ�SP���݉zq���-�-B4��K��<�4[��^ܿy�k�LO��+�K�]�/h)�ke������S����V�m'�Y����9�u��$�u�>ViQ^�B1أ��:"f���b�}T���X��n��lQBk����*���'��]Nq�)V@ƶI��J�$a~�[���rg��9s����N��5��s�k�N5�ِ��E'\:P8LuA˧iw���$��