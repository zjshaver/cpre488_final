XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���G:R���Ql��.4����cD��ޠ{��a��h�eܧ$D�X�tn���M	Z�H�y�Py�ŻQ�i:�K�召P̷������݁���M<�O���)^ۀoU�/G���m��Y�{u�ZO@e�cF�Ǟy�����`l��dcc�>��.�bu���g�!E�ZK/.�z�v��y4��ـ�n����0����|w��t?Y���������N�b���_�A�}�����%��Cv��F)SC"�r׸׮�����b$���>�� �&�ꅇq�ؓ�Oe.	��
S�2��*��@U3� �[O&�*�������A��Mb�w7��6�_����̾b�̈́l٠��UO����v"E�ߓ/����n����(E��^�dHY-z�E�źJ��=��/���aǪ�"�f1Au�U4_$�l��Ӊ�I�W8{����HYB�̄;=A�V>�-1�;+�?���v
)���꾴Z�(�}��jsv�@���{p�Np:��B�U.����#!�-���f�������H x�ff��퇹Ճ��hǝ��W̗U�^tV���\�
[��9�%ڗ���:
��a�%h\�� ��M��O씏�>��"ߍ�rG��Ջdn��o�:����0jf�O��b{����3��H30)��'zs����x�i��]��	�(��Q�T��G`9��,�v>�dz�ɺ�����*���,%��L"�<FRI�͚)N�~�=fp7䎿=JDXlxVHYEB    3a46    1050̗�TabǄ�:o6��{C���d�7� ��`�=Y��/��5,���fl�BkLzp�>n��b
D�ö�ǋ��I]�6w�#n�78���d� `=Is`}�c�hY�0�Ȳ�gQ�sg �9�`�S�W�A�t:�����������O�TO٢�2���R���n�Q�|�jٙ�V����.br}V1Eÿ�ئU�sQ��
('@�r�?��3wK)`��ӿ�h3�ROAS����F\�����`��х�#6l��/���@.sV2�F����8-���֠�b�"��m�)�T�V��Tx�G^=`��uw��_��� �t�.���Y�D�cGޒ�SU�Z�n^�l37��mD�[	�r�����鬴	�	'����¼D��,%l�t�k��S�?T>i,���Nf�;�e�
�0�_s�q�9�|!^ֿ�\�	�<NgH�j�zH������7U��`.5�9ʙg6�3ش�?>B{�}�"�ay��Nv�q��&G��/�uc��1aW�8�= �_����.��}K�s�A�����D��V��'\ۢ4�K�k������E�.j9�rv `����?}dE��	���d �ŌԖ���2Pڋ1�6����}��AZ�-������T��h܄��)	p��vR'�B�+"�������n��|����
��.H��� ��dW�qPukjQ �׾���������dxV�Ql_����
�U�i�Q��3�<Z$n �l�N��۟r7�Qn��C{(�Ź�D��g����1\��<F�t�W���(�v���]��m-�̈́m���^y�aY]:?"o����f�Ww�_r�;���A��
u%���b/�R�'wa?�T#�Sj<	��Ѵ6�þ��#';rٯ�9�����p��Z*�����o+���ق���G�.'n��6��2$~n8)
�;Y��(Ix����a��+.��/�����;���ճ��Xw�lf�,�������� ���Q E��l5��_��*�Ѥ��c�폰9H���1�����{h�#�X��jOr��>!��"��m�&�pq�p�p�ɦK�$8[��[:y�.h2�~�x{�)�}=���<�[Zt�R�����Ȣ�5
�X���c�.h�S䖱��^]���8�f�������m��k�<��x&���8{*diQCu�-ʣ3SV:�RY�hq����t�h������'z���03@Q�m��)�_�fǥX�v�t���=��؟�!�o~��H�=�Ƭ����Q|�ȉ�,������a8�:L����kZӂ��'#3$=�n�8����6�LF����Q|FO����SBȯ�M��@��W5�� }�G�^�m�e��"�X{ZeK�&a~��$�P����eJ�K����y��Ě�%�fM~��F4��O�W���>v/�I�HPp�q�n5:������EM����s̸�o��J�.��:f�q�
/���%��ac<*Z,�r�SH�����G-�Yh��<��W�|���˨g��у�b	6r@�ĜR^vq��c��W-�U�Uu��������d�6(oW��ʺ�5�
d ~�����v�:�/�iq��^D��!~ǁX)/�����/�S�)Q|'�R��>W����{���(v��H��bWsě%��GJ���L5���$�$8����`.H�>:�E|�]\����U�����o������8��[u���᭛�J��>�P�#8~2��$iU�����>F�ߒ3�̌
�p����JӥR��9�e٩���첽d���Q���E��a]�UMYٰj��IF9ҥ�9n���c�f���_�zx�?���'��Ji�)|���_��S��y|�X��]��dYH�X�Q��|�S��n��
���L������d��ˢ�y��%����$@|^�*�V�t\�3�]�!c�j"���mS�X[���Ōt�P�78m��=X �A����U�U����`������!���f���̅���]"�Y�Fh�2&��U�
�I��>��gL���[4�$pY�d�KK�Íp�<�_x���kv�_��+������D5�k��"S\9����e|,������q-�eK���o>��������:�!����
���-{��I�^�8~.�K���ֈ�u�+}	�;ڇ�J��]w#tdݵ̡��2�(S�L{z�u��󠘓II
�#A'.�Rr��fhj�i��<��zV�"�cl�<Ѧ�]U���Y}3j=*��3���ٹ���1��t#anՀ��(k�~Ի\����3������1�p��/��4��R>a�Qd��tU��W#�P��0����r顽!{�@o�;�'��5�h>4es?ˀ���cV��{b�+�!Nc��-0ߕv|��7�W���c����+�2����׾;��6��I���,��걂l�-X�s�0���ݸ��n|�eG��=r2���R�bn+�'s<G]�c��V�ZQ)&�P�L.����D���ا"r��;��)���.�ʪ���4��~�#�m�ޘ_�%l�}O��|�+$�/�[��~����2�2�i��9�/F0�f����e��`w�>��x��4	,L�HvP��)�\i��RMS�x�"Z���'<�������p�\x�/&�1{u���Ȱ�)$�ũbْ��r�@��m�У�`u�s��$m��p9
8p��<�Qj���w]��x`4ꁳ�i~IH� {��`Ea�&[?��Uc>�ՠiV��+i�n�kv��ϕE9�!圇��$� �e�>&��8���%���dH�<�h�|���6V�%M�5�}�)�!�.��בd(��'�Zr
GOj�v1?��洿�*5��D'�lH1�j6��P�u���<�����J��x���u�0|�.��z!2xz�Fi�ʘƾ@ڻ��������26Վ~�؆�/{+%[�m1��N��JcD�:�/ȋ�S]�H	a�)�n!���"�_��L�\bcT�+�zLRO��#{����C�5H�B�#R��� ��:_U�X�[3l
i�Ua��.γ�
$Q��'�i`�m���Kӟd��|�.n\X��(L�֚�P��������p� �q�'"@#�wb뚻KO��jߟ���V7E_d��Pä �(�^�d�����$�i�ۃ'm�+�����X��|ub̹%'���/d���kн^ڄBi_m������M��#�u���*3݈|�,^�[c3�F�Ua���)ԭ��#�-��1��|߶D�@2\󁍴L��͖��ʷS��!1ZiFo\A�˼�P���4��v�I=$��^��Ζ�pqb��HY�#�'��2U2�cZ���/���s�;�l�ڨ$�� �FI������U������1��y��j�b�����W��[l�	�{B�v�Y�*r�gH���޻�Eo{Gf8|T���74J��D�9t核�J�s@�z����Ye~��DPp�[5��)����?W��:d-[<<}��xL�}��[�F-�eJA8z��3G�4�bza����x�B2�B�H�Ӵ^_��~�	[e�	�20����R�x6��
�%S�6X�_����V���S�g�ʾ�4R�U��NN!��iT
�+��jK82pg� P�.�V����M��l*ݝ���6��M8W!�z�G.N]E�Id�~ϖO���M�x�\��aL�#���A�3����%��ɿ���@|waxV��H�DD�f�KGc3�ف EV���r�����B�
�6.ySgJ��ߩ�Z��^O��0�
�V�)K\��t�ݮ&O�����/J"��(���ze%�L(~���FJV�K��9��J��P�Hdɿ��<Ű�B�
3�זU
W��;盼y:��$����4�I�4��dnòQs����ݷ�x��c�W]���������iی�r�����sZ�p23���eZn�(�I ��s=�y����\U�i��7e��ԟ����A�4�m��'1G��Fʛv�Mw�P�$z|9)�F����C7j�j��˼�D5aĳ�o:
�η/�����ɮFø��q闆A��#v��)0p�1o��<�