XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��z������̒H��τ8�I�`d
����u��I {����k�'V缡j�G��;�>�xz�C;Jб[�\'�y^�����z��cdJ@��EG<�O���O��LS��+֐At]�;�+Y�Cvq�R�2��4���L32c ���jy*E9�t�:�GӇ��Ť�K_�Sa����n��wp�k�(S=�b>���w4����t��D�( ����BÎI�q�v�3����Dk�u�k��U�aB+�2Df��7��H���0q$�*��!���^��y��aa�?���_�pV4�RS=�!���i�Ԑ0<B�@
*�[t��V��ċҼhE�IuĖ���\3ue ���dB��V~ ������6�sE8�__�t�)$���ڃ�˱�j�W�hظ�\N���4HU���Ꝅ�`�0)�G3����)gY�x�e�
?1x_1/qG��[ze�P3�Jr�ː2������i��Z:w�1G4o��_ݖP�Oͻ��z�Np���b.��?�ZyM������:A��=�/��Л�Lő�q��+�ۓ��������>���,`ҹ�Bp:�8c<��jn��8�O��T\��*j�I/+�[��Y���AS��*�0Y�������z���a	ח�O?��K��D����nSK�}��RM ���'�C��#	X�?7\�Z��������Хe������6��u^*ٜ[ �w���}X������d=����J�&�mw������:K�x*�ىXlxVHYEB    1a34     990c���C���t��nE��c@�>Q���/�$/��
���3�U��e;�Py�km���}�;�h�����(KTRm���'5�֦�U��4BMa��	��R,�Ӽ�q*�l��_־�A5<҃<W̝5�0�f>p�M��9�^-7��8
�e�"���Z�k���h���8���
�mHJ-+ � �Vo��˽������n�;^}9+ g��d��¬�5J���S]&��P`��CI+�p�$����f2]�ʻ��P��'���{�����B�c��ի����i�6�^���`��I�L����f`d&���a�xHQ�R&1��A�
_"�t�82X&`���'�+_cS���O8�5a����y�Lpq��{��/��K�2��os�B@�>��?,Z� �����]�m��$��W���j��uhשC���E�Z�9��+ޅ���)���Q�ꠡ�eB�i�.?�y����9�J!��,alv@�#���Ñ�s�]��'�ж;�o$���� �ڢ*��ut�!��]$3��y���s�R�.����[o���fx�,ٙ�������j�ĵ��e�Q���iP�}>XH+M֑L��*��n�_4 �F��C��3���r:�6@�\� p�T[-/�H<D��
�y`��6c���E2��j!��'<�t2&�#����Р����9�ɲ�X��/�n̚O���}��,�ۂD<I
h���Ø����;d`�?:�Ʊ ѷ:��r艕ζ���.��v�E�IN�Ҁz*��D�����A{�K���T��r�8����EzDe�}�9v����li�l�NlԵBxbCnU.�oDȄ�c��:� �g�&�km���ra�SQO��y�?!���Q���/�<.�X�U��$*� �g���xW�:/	��V^����[rX�^�m� 瀧��^�m�3��l�n�)jWvr���n�T��p�_H�F^	�Q��,��Q;}Hפ�P�~y���'���7�ѵB?�y��1���&֔����Z�25Yε;su�ԧ; &1�Ri	���=���Z�C[�D�sȆ�h�Ͳ�w,x����V^�ց���vXV�ꁑ����Iz����E��e|��3�;e�x��y�=S����������O��KK� ���4�	I��D��#쌹�V
��p�$R}|Y糸���h���6���W��Pf�(A�m�7��u��F�͸8sPKk��%�=h���9*���JC��=m���(��c,PQ갓r�8㉊��E� �!Зt�����:�kx.���H���ε+���;4���Ѽ�$k8�q��U����J*�(��ޣ��l����m��̾`��*��@�A���x��W!��Bx?�bo��xյ��j��JgJ�<��>N,��3���������2�i���C�r
��l�渥.Y���⫬��B~*��Hҕj��� �g���{�}�4��w�� ���▒C� f���hĥG������}��mC�b�Ry-�,�0$+]>�K,�U��ح|v�"}��pj?�O�ח[K���	�r���a}w\�e�-���5��yPK`��}����i9�J�y�`U��9%n6zׅ@O񙯦�!�ʈ+�2��=�̍�wr%�,�u�E�����`5֋|�~��7��!�B�L�e�$+Fw~������Ui+�Da<K��<�����T���;�o1��n�f�c1���1^�g��t��/2����d��}fc�8NlW�-N/P���1��Ό��bţ3@J[N�o�%�.�ˍ�[�O� ��������Ss�ӳ8g�{{��9�SW��b�� �������d�V�;
ٶ;:�ɡ�]% ��wi�9�~5(!���N�Z��� h��\�=aXj��YH��%;�h�6%@c5�:+��׸?H�G_����.I�����vL�l�\����[;���(�}oK�I�F�_�a��9�K�`%���J��q���,�m�ڵ�@-:�&��5o��w2!��G���R�p<������sm�V���r��~�L������^�-��W���fٗ?<06裱�Pn�썎�p\��}ڢO�N~�Y��.���ɭ�&�Bw]��2Nu����k���4L��|6�ؘ�GI���]K���,�
,����t��y�qS9A�:�.��o���`<xc�a����9�F��	O��9܄�.i�-X���g0f�گHZ$��&�Q9b�(�g.�\�yZ�&f�B�����sp�.�&�+O��;���s<k$YD1�Ȥ&mAI��	��D4��ʒ�w���3߼G!F��zly���x"ō-�܀�QG�>W���Ȟe�+!����M3`��<��1�5|�n/'�ᵠMɺ9