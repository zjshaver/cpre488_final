XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��6�*�3U�	ić�~��Q���ޟu��%�����K>&N��K�ñ��r���^M r�ed����(jb��������{��:�"|���K�i��kl r"��3�?S�ay���5 T��O\$|ŭŗ$�v���,.怸H*�.�a3͠��Lm���"����fI?e�d��)֊+$�E��M�$�	ʔ��=�l�=���"R�5���8SYo��������j ��m�Ӯ������{�=�(����#����9�J3?I�p�Â@|_Xf�tVU��|~�k��s�ON��M��^���7��2��iRg��s�����Rˠ����E��5�Z>�&甘�-�[���gYM�S}m�D��I�sĉCi���-R߀��hc&gW"��c�d`�PH�Z����]pI4��a���s��V|0n@1����p���{R$�T�9�tu���2~5�YqB��L���:J#_N����?'S�`��ލ�����V�y�;*
�XT̅���m�u���Nb� ׳�^D�����i�7�Wb����y�WD~I���=V����63�!
J�Hඟ I7��ح�>0"R����ĳ�/� *�KMg�3��I��D�Z�61v�JH07]�ǫu�G!�G�h���v<ޘ8��Z��12c�p���u�x��)~Ԭ�Q�$�R��KJ���a�(�d�hSƧk�̲������P2���;�>s��B��Ϯې��<�%L���Cv�zXlxVHYEB    374e     ea0�֨lL�e�ېF���;?�"@Ϗqg�|'�JG���b%7Y>�냍�v$�˝u�:�(ttnP���tZ��:���qKE
�۬���*(���Y�ܟ���GFO�~yLZ��c��Vf�1��X����Ʒg���o�6��Al�*c��S�\��O�MA
L�L��+w���[x���F��}����,��C��o�j�����8]m�4�oތ�8J��!��_��h�����V5�P���x�ޣ�݆�/BԐe�����'�`�= �>��m�^52����Od���]jtB�Ɉ������ߌX����^��]�[N݁n~�X/�t�T ��
�����e�j���ea�3zp���i�M:���!�������%�]�$�9٘�¢G��ҁ�~�٠<��C��P�o	��=��dR$bȋ��Y4^�L�'��Z��l4�~��w"�a��+�5%����c���l��}*�b��6��e�up�.]��$�#OE��,L<H��?В���C�z����txS�Q0C�eC�4<�ɂ����.cy�˖�j�G?[�(3�zb��\�R�ф?a�E5Y����o�����X���c71C�x��r�{s�e�e	jcd�
��d��|)^� %�(��3�-�	���|~�a&�q"5�8�g8������~q�QYyGҭ��$N
a3�0
�dj�4�4c��P%��[皹#I{�Ws��a�,0B~I������SM���i�/Ѕ�U�/՟-���[:����uj۩��խ�:�l��I��˟����:���U4�k6�r6i�p<4j;<����c�b4C%;�}dѾr`��S_���o�_OIj]���;ˈ�س	�)&�E�i�E��KRQ��%�@�$j�U�Ȱ1�a�);��.l/!�yP������@���U�ZX�v�@�x���\�=�ǎ�;�i�rrO��zl|u�e�:���<'�s���G.|�|�Z���z{�x�
���D���w�� $f�e%=EI��>�'�#�к�-[^��	:8�ͩ�,�ڌ�^������}3�$�4�A�>-�u�:l#G�H�7z��n�̙n�9�F�oj�&C��(�C�P@�V�����X�ܱ)�m�_N���e��f&���*�B�m8[��[�6�2�o�~�m�}`|Z<H�̡�9O�+��a&�řLh%:aMOb�

+K�(��5��b����>�γΝ!u�i�4����~�ϪP�]z�>j�P��1g�^o��ѽ� �4�D?^
isͿ���3���H'o�l�Ͷ��rې$�w:(������Yg�X#��u�r���]`(�W<�G���%k��p|�9K�R���Wf"��	9��P�3*��Ad�W���A����TX�������U��(-�WAiQ���O-�/ע�ҡ�d���<q&���]A�:N�d��NZ�y �I�����܏d��a��o�̥c1tu~W����P�Ĕ���~���C2.Y�߭��&:�
��*d g�(�"���.C�P�ND����j.�l��H�'�s��ԓQy�摚Yג�4� 11�h=�JqԨ�T*�k�8�J�9+O�|����0Ӯ�}�֩��@:C��	�	�1��ai��[�E��e�5�3�������Gi!��#�_�|/T�{'F��`"�.�~F��H-��G��+�OI+�#r{���F�vf��4���gJ���ꓳ��(��hx#�.W�����[�2F�@���8�S���t'�o��*��j�%Z��'�����9.'���� ��PM`��3��r+���1B(/��y�;��x-�W`v�׿�k<i���VМ����U;H_��$��(�Yoy�I;+6�o��A�	�*��h��E�N�W��7�^�$" ���H��������t�E�Zmݶ�!L�ɷ:~>��\OJ�3�~����A�+�Z.q�B��i��z�٬��]vPQ)(��<G[�m�?�IV��6�S�L�C�[��� /;�3��NQYi�|D�
�	�78�g6ZZ��C��9' ��^�_p!��/�k*��@���V��	RNe>t�It����P��p0D�+w�p��\S 1�M�����a��j�ߕ� <H��Z\s]#���?^4[d��з?[m�s��=�,�C�\#d���WTv�wI:�X�(�E,��`h�ڈ�T�|M4��p~�~��_e�4�.^��:,��5��AK�DX�㫕1�Ծ$=ل�	Px�Z�D_�T�n�D������$v�r��>���rh_�m���ӕ*���䕎��������AFƜ����������J7�l���'�f�-�7���48)�k��r��'R	���wyO
x�����=��VRn�,٬򡁧�B�A���F9�Lw�ҡ�B��sk����� �$t�ۨ�3��!X_���-&�żԻ��0E��k�gz/a�v����QSkAo��������'�%$t@d�xG�̈�.�3E����uq=f�>ѡ+IO(/��J��CZ-!}�*�p�Џ|���;υv�K�t*2��'s]��	�a-��0Xiu���q������C[5�
>��c�jx��1-�7��M�Y��Z�@���]�l��P�F�ǀA;%r�j?z��+�v���(�T���`c��6�5��/���!�2s?1�U�h�A�?����� �ʬ��l�s���Pl75�,����]�q�<��J1Y �z�/|����_x��.�NV,��s�i����ѩ%���׋��]�ӷ�JU�1;�apl<�$���|�Ҿ�B0z����kJ>+@�>B6�4�@��)��&ԩQ�=�����{=�*�����l��IJ�)�y� �i�[�����Y�f��:�-Q�  ���8��iOJ�t|_f�	��u�&�U������L"J�Ay�S_����㤐�S�y�Zq�r-��}YC,���Ҏ���`��%[`4:�.�Y��\���h�)��5ɥ�����̿�����$��~]%��Y�V�x�u�0�Y��#�ޝ���|�^���[V}�~��3���Z�@��獰����g�=����0����ط^���u��Sȹ���i������5��۸�ll�F��o��K~)���t��۶��+����&
 �lLt���ab	0� ��S����"]^���6�>6�6ӎ�N{v0|��_6\m��V��C�<$�}Mlҫ�8��@ž}�q$f��i���vH��:�*��4H��}���#v�Rl0�K�l1�o����]FN�l�Vo5��/p��_:yI��졀� Q\G��G݁0�*�uͲ�����ͯH~\eYI#��t )��[ׇ���9�t�i$3ܓWE�ae˄���f����:�1�D�~0��5G-Pc$R8!�9� �o� ���^牶�2��P��(?�/-l'U1=jl��8Sh��ef&g�>����G�U����&��:�0] �:ɨ0F���-b~�z�D5�^��dV���S���V<@��% ��ӿ�j�(�����2F
ŷdk�x�՜T]�i��;͚j�vb�>���|kh����EY��pA����4K8���2�`���I�j,P�v�tV�bm�j���r4��n�G�(��W���f�