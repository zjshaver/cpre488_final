XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���A���0��7��J�Ġ�m�̐c�q�L�������"=�Y���(�O&�����v���u��-rr�X�]B�������
z��ت%cTr�o& S�?�a@���+�M�#����:��܉���#�B������>JO��/^u���~d�_ci�CA���;�5+x���z�	<�������ZL8r�Ô��Ἰ(�,K��)\F�3P6�c7	_�g�Ja�A�w�����@��?�.�<���j��/^BGm��XK�5�1�|��
��\9��7'
[��p���8N5/�����6�5W %�������A��{��K$������5fP����>���$C���؝�|�[�6�Ȅ���N|�r�2�i��k�������B�x՘��T�f���%��o��Z�B����m�����wA���݂߯��D��$$:F�3/f7rAm^س���vU?�&�B'p^s�J�"o�K�tב�CG�]�>7"�x<�0�-���r�!g�R������ȳ���N@�����7pz�V�"�jqne�9��CS��';q}
��t?	 �rP��|
i�O���-ije)X+R>{m��x�ۚ����q�hݥT���c�b�Ա�{�{#���������<�Ȃ�����`B�<�	Af���.��$�c'
��塌j�~x����/��e�zq[2ͯ�,0��o������B|�[Ot��;�%��bi���D����_�x��tH�XlxVHYEB    3d1e     fa0"��R/а���=:��~,�����Fr�`^��<4�0
R��=����;J�cDHM-�v.)q$e��1$�Z8�z���f��=��2]����]?�sʆ������d�m%���G��5b�#���Q�J���}Ic���>�[�fzwpJ���j�>?���?B�@ Z`�o��lO�cr9{����%��=�TJ�\^��ؙ$��@M��bHpC��ɵ<�r���T�1<����7��QГ�T��_!Z���0$,0 C,2�n+f?�;B{�����m�Q9��g���w���s;��2\y�?� ��G�~�)�G
�<���#/.�Cq	|��ǲ�� Υ�)�`����wS���bcl�"4�t��;��=^�ʞf��%y�
E���!&���_#��-h����i9�l��M�A빀K�b5�Cg��v᫺n<4g��w$֛ �V0c��� Uuv"4�yD+s8��`,l��"q�� Ί%Gi�J�F�eg$jp�����%�q��5���tSK�$�Bد���>����S�N���g+�7��f$.E�R��^�7�?~1ؔ����!
d��Is�]��m�D>j�O�E�0���]�>�pН���O�J@��p%를��࿵)���"&òR����߼$�u��%���w��`|��r�r�x�A��Gcta���Sā���w��#՜�`\2F����ג�M��ǈ �K;<��֢��Q�?C�ı_��xq������=&�ƪ���4�a�_����!�2V�E_zKv�ŝ)tC2X�϶��ĆٓĽ�� ��C;�v�U�ݖ�{�A����I���<<�Q��4�
3i̦%����T
~Ls�ŉ,,7�d����Y��#��8�K���K�'WTp�)�����eq��g�j?�w��a��,^��s�eVF��S^p���9��9QRZ�GS�?�PK���?;b>��x�V��1���T�ԫ�'� �nQC��M�mH����t����5��!�x#^���	�/�y��Y8S�����w�?Uz��â��϶R�<eZ���C�;⭌*��9�'7頄���G�<8�C������*�-�0�����28OX��<����������M&S��9��7ɂϖE3qw���@Ɛ��rW��<�i��x��S�����W�&[�䛼�����j���{m�!{ZC��t�.ʬ�
�T����P��g}Č\w�u�.͍�I��IvUO����8U�N��e4:�� �Zm*��O�ذ;k؝���ٱ��t���R�;��m��g��hNZ?�\"*������ԃkd����5s�����`���>�c]}C��U(��ul*!�b��0�����r�!.��{�pt]�[��-��� ��?�"V���Θ1��ۄ�gW��6�/9�G�Q�&O�hv�y�������O�q�\�3�h�܅��p�?�+&�d)-��Y!�S׮���}�9��	E:B0��VPA� �
�+�)7�:Ό� _�{%��0(9��n�Nk0p�"F�5jR�u��/�P�^;����l�N_�/��#���V�ݾIO�X4���_�͵!��T�h�zV���=9�*:\�]��F��~�i>�Uf =�0j�����x�."5�8�°�:l�5�vD�)�|�ƞ�Kx`%+�
+lGax��7.�C�)�LX�i�&���Y6���` ,����C� �q���c��S�ĥng�|{�fm~�4O���82���~&�;�b��l�1�ߏ3#	*�.4(�P�n�~�,c����x�5��6����z��oe��:��VJڪ&a���7W�桄b�P�)`��ڹ�$Ѣ���8�/�FL恧-k��>��ZhyF����$�9�Vt����"�dD�9�<��ܢ1�Uq���Ϯ�	�������E}��"�R�P<��m��hQ���MA,H���Rf�sK��i�ʍ�eV�S6Zw��:ys�E]#��On64r�b��<��[�`��"�z5!wj�!xħ�'X�s�*V��<_oq�\�-����N-�,c���'���a�Ce��/51<i�]䠊ܸzZ�DЮ�TD�q�}Gx6���=>��sÖ�_�Тx��t��d̟OOW��BҒ{U�`�s���yfg4�.ֺ���l�4��3�F�֯b����a ��io��cA��b�0��ö�k*����e�~t7,٥_���t⨏-��1AP{gF��C�;
���TE�*�:'0��O�B����\���ͨ������ ل����Q���\
��g�fu���4����,Yo�nQ݉��rG����o���#��5�.����rd<Jև�'��zߛ�p>�.z�@�(u+�S��<��oR���|&�M�>7�#�M��Ύz^���������%���
)Ä��� 6��ǫ�9�R�-��R�5�GA��l�YS�_��~U������1����-�v�;�n�ﯪ���4�`ec��?��AW����v_��V@����e���{f�� 86A7���>���O���r\Ah�pK��w#�	���{���������6��eK:��2�y��<�5ȉ0LVmҁTl+����?�x�5�_�	��e��DL5f����j�>Z�`�����d@�(��4�A�)e9dk^ @Y6Y��"��� �Ľ������2���_�:�K���i��g��o�#,6�̴�~R�-:�@�H����x2�B�'q����ߍ2�63��F�}~=���g:�b:����)����ήxy��.5�$�-�+�ۄ���<j>��W���iB�H"�w�7�eM�u5_�����}(��؇�q�2팜T-K�E�w�2Zo�I���W�
�t�cQ�	�&ȾOd;����A��h�z�Ѳ𜊪�0;ؔ�B�ʕ����H�l���O����#]�,�
���q����Paմ��6�SrFa
�<T"������evQ����ZSPy$Vv�g����"� ��3�X���
�N�d�?t-��l����\���"k��# �5�C9�<N�9�vo:�9<xU�)j�������${S�G��M��U�.^#���łb>]؝f�O�#R����"#����o��;�y���zZ�+}H[F�p6Rp�>�!]��G�M2��T �,����x=�f�EP��Kh9VF�U��9���#=I�u�:3-ޖ�|��hL�Y�d����/��y�)uŉ� ��
�4���yBw�h�;�%���*&��\,�Y=^�o�����dwhԲ���n܋�N��S{��ޭ��ܥG�6�|�!�Om_y�^��������HJ)��*r�X�?[�l�Y�T�Mo�q�m��*�7��&���O��±��8{�3J�n�갭���Ɏ^h
n���N;$��V�Z�r��;2J�H�~���/�\������uRjl=�4u9CRM�2��e�n����ۧ��o��v�
�o�B�nS�$xq��"�Y��)Ԍ��w��9�/��rS9��v�cBUl�nmP�zHg���/��	�!��=%��c�zᡝ�xb����;��F��W�����}���:1)�����X˥$�L��s�t݋HږQfR�Ǻȕ$�.�S/�!>=��-O{9�I{e
V�� [�'}�<�*��Coew5Ċ��)�J�5�_)��<���C���@�Þ�X+TnL�r�&YHT��,�H)-z�턃J��q�H�ۦg0�3� �Rd���ժ�1X�����;E+�+��- �~�%��H	�_����G`�X�	�Ox_�,�/L���g�^��)�԰���u|�)�|hz���[F����H�Ȗ�����=�S�Њ�mQK�o�>�m���	����_~:�)V�j