XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��.�.c`���3�f�|r-���s�E����k%r]X�Z�dop�t(��b��?�b?4�͐<!����t�/m4�V��z<ќ��|v�����X�$l���Y!�<E2P�}�.��K5D�{ԇ���su~��=0�m�E�ӑ�p�����`��$r��Ї�MC�(d�0����Ӷ6 =^G��i_��g��A`�cN��(�2s'J�W������\�WzrRzqU�-��я):XP��7�!J�v3j�]�{\ 	ꁭ�8//·�	9����֯��(��R��]���4�C�4נދ�MH��8�y�HM�P�H��=*��s�P� ��[@�{ϒ�Ѽ%VL󣨗[߻�fX�HZOn��
σJ��l&���Kd��
u�S��d����V�8Mӵ�FGo�w"&ZY�F��ֵ*0����^+p~Kݘ�?�G�A�J�{��sn#N.q�j,I��ֿ݊i^(�d|����u���&nFЃ)x��\;+tʥQzu%Ÿ&c�+��ls�ڋ!���@���O�:}Wib�T��U�3�i�QX�-؂��4|�60��3i���(�j���;Cއ��8�Rm4�&���9��-���D��_+���ѱ��3�1Lz�jY_֙iJ�C�mѹ�;i
��|dL��QN�4`l#:�l2	�#�}�P$.<�CXy�\��z`�g�5J��ZP��1Udl��"sO�֯���9R���jb��h�0�=tW#Ë�7�y�F�pXlxVHYEB    5d29    1390&DwO���|}.��Թ��«ݰ���.��BsG��Ёe����C�.��4�g6`F|�V$��rH���w$I���b���^î.ҽ����b�{_E45֝3�v}K��7�����F9ڮ�p��6�G�vC���UڛM B������
�b���-��m���]��܃�,Fm�%) �Я�0a05��	�0�G�������V��?	P)2��y�,Vp3Ȥ���@��.�����XM�7��'���Ɛ��J��;����p�^�����f/~|��%�(�20���k>���G��:���]^[?�[=�j��
p�I�؞�哺�N�P�i
U�M&�3��lye��}t��.���,z�:z�{'bwߓ��X�+nBV~W�v8�c���e�6��F�a{�Ճ��5(�F�����|o)�A��ód��.�]|������u�@f'e�]����!T�=���Z�w�`2[�c�JKW��lu�a+�b)Ǟ*� ��kI�A
Ѳ2q�u��(?����P���W�M���ň'Ç�3S������-�yo=�7l�0]Yؔ����mE����|�Y$��}�)�t����wZ �S�ȃE�İB���y���ޥ�:ߏ� #�j��CY��WO&jI5�
%(ƻ�Ҭ,c�h~9�h��t�.�/V
��c��+�?�F��'��Ҥ��Χ
�<ب`�A�I��c��7�@�=J<�[#d�P��ްE�u��OF]k�������@ࣂ�����`d�4�䞐*g��`������g�X�?Abzx2Dԑ�֪�md����"a���\�z�����"n��A �p���7�Wb����Mw��Mq{g��z��˛)�R����3�K^�P�h2*_��{�2�5Mr�V���ty��\#����A��N��n�"�!����K3��|O�+@�k���aF�{��	��Wı���e)P��_�M-�_T�Ȩ����vY����z����g��Ä6����Z�!ƴP��1�%�M��v����қ�&7���Ha�]�E#Ga��?��~����b�j�w�l&��sxEKc�M��VOd�B�y��E�ק�:Z��0`���� @�om�'9�rT�%Y�|K�Kꐳ!�W�~+����Sg�Cod7Z���B̔R��E�+ظ�!��x���z�[�="%���Tg�r p#Rt,�>�}�+PQn�ƾ���D��'7�; 1�e��ȺBa���`'���&������i�a�: +Υ-ٵړa@��K'�^�12���P�Y}�"��A�dB���:��Σ�n}Z��,j��ܥ��)Ԫ�#/H��睼�7�[#���"8�#��>=���B����q:����H
����V�H*�gǥ�m�M�l����'֐������ě�!��{ǐ�U�|���Xg��1��7�zpO��KXN��r��"��e�ܗ�R`Pkv�f�,'0YA� �#a��>h��^A.��[ ���CW"	�N��rT�I�n�ԗb�"�$�<�0���n��l�;� �l��j̊�	�y�6�������t���&�K�{�y�f�ԣv6��q�� g���f��oP+?r��<��lM��S�\�3�r~��V�8�L�,��OAx߹�1��(�Mvx8�6�3�e����E���a����KN��hF`���h��$c]�~��i+!�ak��-$]nG%=ڢm�8W����%�!,�3��C���s_v�B���� %�(��Z�Y� a���8h�/�J� �wm����>"&^Ȝ!H�Q��1�����w���[��HV��[���i'�0��LCKmJ|�Ln&�)��[1g��M`+�{3��6��h�M[��u��V��H}�����F�J�_���O�e���e��gGެ���w�/NT�2F(���X��	�]Ci6~�=�,��e˂Md]��U�v�ԯ�2�lxώ�������=���v:�̿��F����S8��#������ɱ0Y���)�E>�:�k�!���i�zJ_qM0�U���]���s[����Q�2?�r%���z�S���cd�d���ED	��`X�q\;ULOKh�/4�R�Z��+�e�{��F�,�F4U�M�R���u�I�D�����'��6pG�z�$4*��L]BG�6��#�	�|�鼺$���8��m�zH�l�va�p�=G,�-�H��ȼdN�>5g�By:^7����hB� �6�]��c�{Ή^�od�� e"f����n��O�)�����	��E���**��'0�mu�ocT�r�#�g��I���D�|(���{@;�s�$�m���%���f�>V��a�Q�$�l/������m�n�83~]	�(�ߞ-UA�9Ky�.�Fbg1��ٴ�Jy�A�
1t__�ˋ]�k͉������`�I8��-5��TP��ο<�3H��|V�?����h�*7�[����`\+��w�jQ�$ث�2�d�s�p��C�le!{�٭S���m����`'f��s�}D�J/�
���:��X���ݒp���d�i1}�o�T� ��._��nVD;��:Ql�i{��@_9)��]	�����2�a�c��>l����3��M'U�D�1Y�4�ǰ����[�Րu��5�'C���)u�*Uc�fB�9�7z$i�~���>`���z�t��=5��|(�:�h9(ϪJ�
�|ˊv>�s��l'
����/ЎdZ��|G�ag��MCYZB���r��\�ճP�8�'@��g��Nh��e���J�|c�(L�ueS=9q�S�ߛo�EX�����k����^��z��粐LR�&��� h�x��/�_��\�ݢ������#m�T�������B��yݡ|��z�����;pSҔNL��E�#����l�a�2N����N�z��@��e�8Fэ{\Y	�e�XµVH۶dܠ���BB�@�t���t�f$]���
qLez6��6Qc�NQN�*V��&��|>� �2ZϺ(R���b��s��Ί4Cy+���ٱ�]��,6��6��*��	[�k5?�s��s���J3�U��t���� w��*��sO����z����/4�3:�U&x��P�o�k��@p���Y}�:��*�XMG�ZvUX�'�M���I|��?�4�����#� b<��&H�����!&���KW?��9,�S������	���[}5�h�5�n*�!�_~@�2�`ⵯ�j�����`��o˃NC�����$U 4Y�'4����3f`�?��8dPg��*�Sm{u��5�� �$��	?!MT��Ь� 0\U�Lj�As���T�7)���az�x��:=��ޮ8ԏM٠�702�Kk�Q&2�G`��	`|���I[�����N+��8�����������VGLW�E���������Ї�B��lB������/��*�i��q�
��6����$aj?����X�|�5�=黧u�}�x��K��z ��\�mP 2vH��I����]���u�J$����B�-^����L���T��LV�dB�����7��&L��"_oPp  �3��������(�Sy�&u����L��^(ۄ���j���!_���qJ�b0ʷ�t���:��$e1�Ӑ�l������GE��v���M/�>��̈����z�$�a�P��Q�ۏ4���K��>$����l� v'�;�Q%V36\:Tv���H+f\uҡ��=��~��.�K�g�:���R"���V�U���(��k�Q�#�j<9�x�1s��-�_��|j���}��=�D�Ԇ�A��Q��[��x��en�q�Kj�W_�_!���)"�m��F��U[��ѶÒ;����`W������C��0�8�k/�uU7h���*Q�i�E��^�Ύ��Y`��u�[x�k��ԙ�)sHHyt�����*�7`b�d��>Q�_0��	�q<���1o�_��ٺL��.z~�/G��*���P�ov�#�؏Ofȭ|3��'��8~��t�� ��5�7��2`�����\5��Ua6�3� ;��lv�>(ߋ<�*)���M>��{���$�������Y�Am;�o�5�#��ж��j���t��>g2&D��j��b�3���4��Af�]M�<}��E���I-�	xE�����ό8�f�y����w�ڈ�d���p�|�Pyh�ݤl�.�?��6Vbl,��>C�S����v����|�1�y� TnT�"��@1�N{
����e��s��1q#K0~1hM��Je�����������S,A�EI
.�<rS���d3�'{nU�_�r*M��o�T���bj�F"on q�؆ī����"�֏��+��R�{�r���g�|d/��!Q��%\.o�b�%����QA\Ȃb������y���.�'�i�Uۆ�(�4��_K
���X����� az�I�w���_)"��~0]�8�"�y���o�	���[& ��gup��,RH2e�c�N����ʣ�b������n�?�ǅ9�r���m���+
hrg�����I4���0���凉/�z���p�Y��f��J�����gy�2�.Z|�0B7��Ч���ܟ�����i�DQ��*��om��,��T��U& 8N$�I[���v���1��ˌ�V����\��_aXs���!�4��߰�}�|������e�[V$�DϿB�*�'p#�G��\����{2qf����ǂ������1Q� pA�Vp�5C�a��f��^6d�x^I��R.�5	<����x��A/k�㖞 ��qX�%٪���H�$��m�.q9�w)|GF*��q��� +il��p�m�co����R�(q�2����,UTe0��V��M#�Mj�X!��g��PFf#Ly1�vk�X�m	R�ef5{{e�