XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��$��O����e���h��IT-Wj�|�d�T�-v:��+M���F�A/�Bv��j������dl��~p�q�0Z"#���ΣV
��%)�D�u_�N�DO�T�hodeS;a�|m���$E���Y~��߃f���usS�	Dq#�Dl��t0�l�\h�2�U��3B�!W�Icp^�c5�̅-(n�����f�uԽU�(hZ�.��{o%2�r�L��P����-L�%y�$*�ʠ�=�+!����(޵��l>h&�t|��ގ��z�
�O1di����>��TTX���2�90��M�� <��yt�n��-�N3��e�nN����u/��	'��/��Hf!yB����x��K*�J��r{}�����E���|���c��Q�HHS4��U����Wc��*�j��)�\�N��_���C�}Z�"3@m�0���@��I'�ά�=���pr��~���C��R��W�� 傀���jCp[q���t"zW�uP��`�B�B#.U��v@C�����ʜ2w�P�z�69s����8�+�(����`\�l9_˩���e�wj� B�w���:��޼7�D�^�	�[8����������d�z��|+�[]�$�`õ���mV때)�lGC��]�Y�)�m`��?�!RV�䒣&UNaY祋(�kg�xGo��I�|P�����Rp�2�oh��~}�؋��߲���iX�+k9��#�]t?E��Jfeht���lQ�]S#F�ڣ0�j	��MZߦ���[�XlxVHYEB    28ae     b60}��2��b��1���N9����ª`[d��x���I�&�Ϙ'm��}���"�PAu��c���!���-K�'v����rG3:H"<��̵@ 2��o�!��9���1_����^���I_p�����^:��X.��*�
��SSG0�?���(�����8�V��{�)6�
�`Ҵ|�$�N����#:yeh]m�c(�e��>leHr�5ڢ($�~�m�m#�k~&wK����E5��\���b�g�9B�9�s�CGADI�<,���u��f��;;�DHˏ�ԑvfrƬL̙)%�-������{�S���:��e��"��x�v�Yd/��UޞB�9����wag{�6�ZMX#K�R�r�=�S��ϝ�/x�V?Hav�)�Ei��4&��9����{��6�S^��C��iQ)~([E'�*�5����.�'���#�  ��pf��L�*�H��&�^YSg�īNT�Ql�O���.� �G�ש'i�{�a?�*�JJ��k�O�C���5AD�5�Q���֜Q94�c�L�ꄁ�b�yAU�
l�p��<���:���e�T���*�W���UA2��cd�� ��v&��������҅��.X����������dإ�s��qnb%� ڈ��8�:�;q�C����~I���.�p��;]�TkVV�@���Ȇ�����8!>�FՐ��_��y�ʃ׬�� ���F�K�5��j��>V1�~e����W�I��jhCAkgV�r(����ڑ��</6�(�6�V��䖝�a�����á
{�G2�Z(M�����vٚ֐^p��K�Dm3@���t�h�����t������q������C��j��?��{�/�y]����O����_��%�U��G��ߧ�.$[J��O��w8�v����+�N�$U����Ie��U�]�%��b@7��Q"�x7+b�E*a���k\Ai�6�j�m42��*�� �#|n�J�CD�ӹ�za[�Z�<$pH����>��n�u��)g7_$H��_󎴹h+��I+�ޙY1�$M��?����$4�C�&L�%wv���{ a��ֺ�6pl=���Ok��S���0���	Òc�G�f�]������ɼc�m~\�����L��&m]Q����%��SB�1�|��Ē���#��x��%Y;�[�E����@��k��F��ZT�f����K���-�_�$�ń=�����T�����W$D�⦍V-�봊����� ���;�'�I�0 L�� ���	��3�]��h�#e���0�}���"8�j���,|:�9�^v������cQ��Ĳ;TV �i�S����G��a�Y�R#kT8=D��]�!��
V�hj%���֎��Y>��#��M��h�a�l�<�=T�w`������<=lC�ݰ����"��~�Ȯ���m��'=�l�3On7����/H'j�b	�f�����%�W���F@-�a�;(��gU�����]�-�Q�i��'���h���e~Kw�x���,>�?�<�P�(�æM��S�!{Ј�8�y7�q��?�It�ub+���������~w�2F�BUoz�uf�a��4}�L~!5�/"���T<�5>��$*�2�+�h8��>JУ��=� cW�<U�D�=������+L��R�OV |�7W�VK��/��2 _>4�����������U�٪����)�?dă1�q�NyADu?��i�PJ�˓�xwn���6�r�鯻��z&���5'��p$�D���	<�A��v�N�uG�%JWk15C`x�>�@�Mc���][��ڽ&%�o��-sI�E�\���'�a,�EM�\�M���%b�wIE�����cժ��l`"�<5�!w�J�F����92a�<j�?��04�Vw������<�N�ђ�� �GWPg&�~{7��tX�;3\{B�dz.X__����Z7z��`n��s���T[��vm�#���W�ߝq!9X�-YƯ��qpQ(�J~L�	��,}�K��07d�i
Q�T�>.$TR����

.�0g�ɼ��d�ջ��x^:�@8O�E`�@ś	)��@��`�b�S����ʠ/�H�?��#`�G�f�}����C�8�
Mfl'�xc���n���j�*�2�egv�3���g,������N8�dM�fb��l����L��x��L���YOtH�*�#n�ߞ�mL�V����b]���?���b�����7��|!LGŽM�q���[0�	aK���;ܐ�l��A�R�jp���7��ɹ*.�jLb��5��TK���ն�T�O�\�pZM����JL
d9!�]$g ��x�M�?��� Xb�W��S�$��u
b�n~�{ǫjd��������=��X��hrÑ�VQN%E�v� �����G�svAI�B�9b%S��؁Hn��[|/Q��3V(|2ǫ�vA}}`H��u��NV�o�dŃ�+��&��z���k��/8���ã����;�_Rv���W�ފ.0��;0C��(0@��eb�Z�'i/}C�)@e=za�����} ���- h���H��:{D�����k!�!F�f$������*��%�6ޑJرm���,�)��4�����	�J��)
_o��«S�"yIHޒ�*��HN*�����v�3���RV�('%K4�ѫ�+ ���_�x.l5}����e��p���b�Eb���v��"���H]�{ZTsƬj7:4Ƚ�P��#��z�{ˊ��P|�/ �zr����`�������FJ������c����֭Y�� �36�Oʫ��RǦ.c(o\"<3-L�Џ��9�	
@�wYR����a����q�D�r�x��ڻI�QU