XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��NSl��o�5��A��6���Cc��˒���0��I.���=CD�.m�:Ծ�&���b2۾a�g�]W
vDe%ղ�trGZ��$�]�5��+��u
;C�S��9+0r���"k�XlĬDda�Y鳄A�j2����Zv\��v�F
#�/Ӆ��ߖ�ێ���02 �[�]���Ra�	�2�W�#��dS��Z�)����!�S\�m!RT%� ���ߏ��Ae���$�7���)� ��{��:�$�<����x�!y���d��
�8y6Rsa���&墏�{�sCr-��9��9�ۛU��H��q傯:}���%yj�*7��(�6��A4ʃJ�RV,�L�lܴ�qmхni�%�`���)�������8Z^���U��������E�(cmV6��?��/_z_�J��"���d-	r���=�V� �m��-�
�}�{�0��'e6�1L1z�#��.��ۄ�6y$��Omұ���@��R���ϻ�@��z��ɝ�|�[�N�_b��lq��>�\o���q�v�.�,���4>6��a��/%j���>dY�{�2bߤ�����c�G�r#d�b���9�Z����IeɼZ��i~.-9��e��js����N��k�˯E�Ht�<�b�#�N��@�A�_^�Y�{�{���T�m�Ԝ$���u��pۄ���d���[,�� �}o�/�cE�M�)�g��Z�ʝ2�n~�nK���$;M�v_p=8{�X�Q��^c�C �hcXlxVHYEB    5e2b    1530>�?���a��R�b� 9�p�]P��\$rN0�s��h�j�m1�J��f����Vq���V�/�I=Y |NaN;��M�&Qrs����z���a���O���HI�G<RcH#��/�L�)A�3��?n�y�X�R'�$���x^م%��gPq��Kp�Q�{�`�"����{����_�B!Ŀ@y}��30i9D�/WC��%��7���>LU�T��i�	�����^{���ɦ�s4��(W�Vt�Ɯ~N�@��m�O�����i�F>�?gǃ�.<O��d7���e��_��r�}.Ml�s'���7i���x�,�O�{s��Ӣ�7k���H��P���>-Y'-���`�?d�^����{�:�����Rf?;� ��s�˪���t��O`��.�\��c�*u�MA@�<ݑ�]!�M��jm�ѪQ��_���i�2�y)�b�]|o:kbDǼ�YU������V�X�#�ߺ�٠��K�{J�r����F�,#�o��<�q=��������Y�Z�X�g�M)�f[��p��^Unе��k��<� C0��.��e�.Cm�Q]�+��q�[�	��mS�-��_�5�������Xν������/����ʟ"8��tǓ�MJ���� {��N�(�����'T��G��8f������n^��`Z��|J���'�t>��}u�CY�]�����qXS�ni�8x������6f����F�[Pݥ)U�����M(f�N/v���^@�WCa]�%2��?~�8�A�����o5�2�5��{��>n4��Y��V��2.P��d>�Bw��ue����t�O��R7v6��C6� �/�i����C�]�]�/����:�jB�{�w2�"���_����|,�=DCj�L`+�H�cDD��X\S��"��f�,����§=X��,�;��+2�=�"�?�H�����C���y���,�x ]��q�0��BS�_�s���,$3�!S ��#+���=������0�.9Px�fe��-�o�_d8�_E�m0�nMr�!��9�]|�A�l�z��B{�'@�y�������E.#�be�X'{z�Q�w/d0(

b�h�ԡ��t�2"UO�"������T[3�\�`N�h�^E?���a����
�~^FT�8��P��~:��K�qfh�I��d����"d���TLY��V��5A���4�SXWk�aBQ<��#Q{f���~�1{Þq�J8N�:���y���ư�͸^�f������=��?�dspRPQ��dZk��l�w\�7'�f{Z)T*s�Z�v�vs��d�♆������tޕćs�Ro�>��a^'�w��~�*PT�;\y��S��>�*h������"O��Z��ۑPrG�y3��s�A�)�X)"�}�`�1��ܞZ[��+Y{I�v�[B�D����[���X�=�E��?#pG�A8���R�X:��:�ɱ"ʺ�$V�hl���
g�y&qȖ3��˥��N���G4��D��{)M���b�smh��E�2ㄽ=�%v,lx\ ���!U��鄾,����
�D8�f6�$K�� ��U�R��?=0�}^�`��ۏ���ͅĴ>������{������|�E��F&n=�ֱ%��������#l�l��SW��u�v��p��ғ���qq����(�FH{ � �p7	D�&���p��ʧ�:��a���*���[���邖��G�l��-��ȶ��b�.����{��+|�2�E>pҕ;�_{��G�H	�*��P�hSu6U���j18�
���/�����"�S�6I����F6K���5+sE=m?�V������y�����F>�;�ө��d�r��x�I�xL�GeT�~_K������F�|��f����"��$B�l*�jl=v��wg	�[Q�s������@�,	�V�n��3=[W�Yf�1�L����퐻>'hf��)'��y�U�kU��9-]2}�Ǿ�(),��Y��}i��jyL�`h�<��Y��V�N�
���l3!|�qaw��ʈ�9mA�`z��;�0���ܔ�9����ӷ���+_[�8���@t (�Pnn�{�'�O�=��%r��%p�8������f�ّ����q�G/*!"&|��m�#���7@�i��>ں5�v�
�xEi)��]1�g�.y3��W_����OK��/�C�do I��`�k��s"���xw��(���|��>��z^5�y΃K�.MZοe ��fS>S��mm��=E��ǫ�?a��B3 8�0o�*TW�h�ݒ�'��9���J�z�qq�F�u~�T�vq��0��h�0�E��w��98�2J8lҷZ&��~�~�?MD�{ �K9o62�n�gf}i�q�+��Y�SՓ�ƕ���	p�	���ָ`�7�V�QX��[6�K����R�\�2��T[�kLHe��/F&C3��;�JR(�,f�����c�&0��B5��5����Fx ε���Bm�|��R�w=l.r��9���ٱ��$u����Kv��(nN���_;E�GA2&1÷_L�'Te;�h�@�S}ރV(Sq�G�ٷ,��41���ڍ<g���� 9�f�־mr�ei�f�)��iJ�v���L�*��)k0e�	#h+~8�Q�@���`@I��P�Jpx���ݑ0�fx�PN2L����w�h��b����r�T.�z"�_��a�u<��X1L�´ۇ۲��  v_��?���=�$��X���_�4������>�V�,1�n���=�>*O��u̐`G���p���@�ϗ��KoF)��"���ר�1Ǫ�_(@q
pH ���zW�����۬<Qv�d����x��Q�B#�WS���g�A��k�:{4�����i��ژ�*�x�K���3�n^6e]����5�.���|[����l:j�r0^$����m���qt�P��"F+�� �����cOO������dK�^�b'��%��ɞZ~\�Q�/r ^h�m��֝�;�+Fs�iѹ�-F�Z�}�  ��G�'7*���KF"���r`ض��A\
��HS��<�VZ������fv�s��XP�{�Qj�ky'��#$����(t9���sM)�,���ţ�}��9T��7{�(�+yX���ےO_�����ζK�]/�B�Y;�6�H˾=V,>e-�K7���Q�d)����)�+��"�hǚi+ j���,�����J�{�4��
}LHF��
�8��Sk�+�S��
��F6��Q���n�5�xg�j�ΦS�[Լ�Ui�]���S*��W^; ?Jx���7|<�j�[��Hb�åW�DY���Ț���=��#�={��H@�ӹ�YeR�s�&Q���'�b���=�n�yRO��}��btu��3¿#(�j~?t!U������(�X���F�fCv�d&�K]f�|C��C�0d�ƈ�C�$��#�=��!X~�}�Y��G���}w���6�h.�.��׍D��N��z7U��օ�y:�P�=��':1�K�jq�!/!�j�]�	m��f[�*�;��Zhv�Z{�"��p�����(�<�J�/���Z�C�|�s��.���NJX⋇^S�v#�>P[/�G��背��X����-�.�0�"�L�i���X{V�Q�L�.�~��%cJ㫊��{E��Xf��Xbޮ�,1Y�-�4uq��w�'���U���z�t��s�����o,I]?r��J�K�����B:�5b�h��qq=������1K���8�&�>e9��q���~�EB����0~�B@x�âx�^��7̨^ʓ���U��op�o�zzĚ���V�]yoZ�,`. y��>I����@���e�K4���Ș�8�	U���z�d�n���YT]���4�N>����V�pTR�O#�^�֖�Ƣ��`0�R�Tǅ%��n|��t-�؄��;k�wxD~�+����~AGw�@B��)�l�%��O��ǀK�pt��8�Ki}����	����Q6�������:��L�#��v&�?�iˋ/H����)o?� ǡ!&�����"]�1t�*�;��)~�������t�'�QO���2\�ϭl��i��jh��ԛ�E	]���r[]j{祶,�\1�-�徍1Z��=J@������KP������Ad˒iXQ��O'<�s	��Qv��Ż1�5 o���w�E���������#�٣��W������O�u�zc�9�"�G�3��k�Bqm�u'nW1q������O��Uŗ�9���$@�,�ɘ�q �.�UǊ��}{A34^y��q9�}������pR�l f<�о~�4�;�|�$��4�J�R߆�,����ɏ@��7��?�v9��+/���!�$�@Fど�;�E��d�nBC!��q�nȞ9t���_1��HX�4^�9���<Ǿ��m4���6�[����4-�y�B����¢�g݋Y��c"&J/��w�
��M6$���YbcȾ�{,�o�b���Ha������)�=�‣��D��܊�d^*�Tq=%z�Fr\#�{��'L����^d�����OM�b-SY�,z�U�,z:}~_�����s�؇�2��]"���SF�kWJi��S6�U_�K��񁦛ǃ�>����R�ėv���j�8����a��WiO+靫�������E����Y)���+;�b��Hy�~��BҒ	�8�x���+ā0s�G:(��D$,�?ih��YÅ'æ1�߮3��_q����~�h�����sf7Ձ�6�)Q7����)�����"�%��-�wfN��3�	-�k���ٲ��!��Z�t�ˉ�h͔������pf�U�����b<�iȒ+;�}��gO�)bp���d�̜����UP�kЉ�&<j2n�"ɂ�����3ń��L	�O�
�K���p2҈f1���iC<��!��cD�P"W=;a36��I�
�@�[�8>����v����&b��u�Y�-��?g��ϢI����SG��t�Ԉ�N
��za¢s�Kt�ToI/w��JʍBb;8RM)���q���ݚz����C��g�A�&Yd�	]o�]Ɛ���g�RC:ϐ�⯮������6,��
��� �^��gs�xgq���3�2� �l������G0D5q9a<Y�A��:X,J �(�Q�u�O��c�*<׫�e)sc0s�
6�R�0 F�iv�[� ��ڱ0�۞u�q�1�}\ZZI��C7A�7����8"�Q�p*p�1�uGj�UY��l=��4�ׇLz����H�9