XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����yr"��3�󬘎`�Fj\/��G����{�->S��p�-����OVe�c��_@���B�/����� R�O*eE��)ٲ����E�ك0�s1��8t8���ݮ�ғ���>���[�p�E� ��f�b���K'ƀ��`�Zz��IY�+<���e�����i��d u�l٦Q�=vw�9��u�Ut���q]�HO��"���๤�T)�.�w�nP��fF���M]�8FY�l��t���R��wh]�������T�G&Ogb��u ��k�q:�E��M͟��\^�2 ��=��t)i��N:.Gu'߸����ޔ���4������dw&��y����9��'���t����u���%F�h�E$ Y��6Q{7R|��~�e���B䚖��$X�:y��	�IQ���ZP���/&O[�M`����qY4���v4#�����_�G|�Q������y�OųL�B��ݚ+�]/�Q�cH�c���А���{����XU�5sm���ZU�Td�c< ��fZ.o�I$7u�����*a՘�3�wtC���7����&�~�w�A���add��,E���
�g�Jk�g��L����ߎb4ˑ9߮��?gVF�2�P`w��ӝ�3d��2"Ś�NqV�Qhq: �@����O|���~yvǧ=�0f´H!5'S�#S8DX�-�4�%�8Y�o�����b�7���0�:�5�M���m���ۡq�8w)a)��Қ�˼�(XlxVHYEB    5cad     f00����^������/A�K<�E�>,5D5�@�S��O�k��&���E	�����M1EP�n그���j|3��eɎl���x/5 �)-��kTp��˻�����H|U���'8�Jj�F��L��N���
�ɚ�Iy��(�,�U��m[�UP~l�sƱ+1�[�Y����N���,�_,Sz_S�<-�O�)�n[��W�B��,xe�š�y�ǝm�#��P_N�"N�~�%��ѳ�����c�0R�n�\�#M��_w��6���}\d�8�pP'����ã�J�)�k.��������
����7#%ȿ�E�7���%
�7�)�;��NL�X �x.�t�y�)������'��C�b�%?l�i����O���"�Ѭ�n�P�H;�< �p\�ޫ� @F+q�p&�"Akǚʙ�ˁ�<^lľZ���1̱����̔%���0Hq��l��B�9��]��$��}բh:tt8�ޙ{��U�A
s��%�p�����Z�h�e�'V�6e�V%��)	�%;~l��i"'d�h�H���[l(��s�Z��ǜ�pﱨAӽ�ż���.��@P�ھ�I�-���H�&��X�lx�"���~�����Q��`�?��l_�f��`Ff&�W�K}]�/���1-�2[���o��Q��.�Qk��f���t���3F��c�]�~�"ٕ5�*��Tڿ�ƃ�BE֑ �����('|&o��e�a����Yd^u��;)�8 �>h��b��_�cTF�[s_1J ���^���#Zns-b3����k���vH{.ץ{���F�v��M9��|�5������B��&��h:��U�uk�:��3��q�>�8�Q�8F?t���Ic�w]����x1*�Dh\��ct ���\W�s�Չз[��u��J�Y4R:R=<Q��������]�`��Ŗp ��(<!��E�4<�Fz�WٻQ^`�Bm�[�c 	��f�����K�|�NCA�ri<!ҊND-����5����i��>�9M�J?���hз�H[��	�ҧ ؀N4��~�E�J��c!������d��+2���kK�I�T�/T��w���)��b����:�F4u�y���8�`�[/��~����s����ve�tdA��'�����?]�̟.+� �p�E+s�,��4�(�U�jr��&��c��1��ipT�yo��<	�t�-:�$��N�U]��D��=d�c���41V��6�z��_��=�)�z>bGO�r2_��1��rH��r{��Pȭ�Td���7Up�kc���%��\!A��y`�c���y���1���\f9�S5O}�jb�1���[���f�R�=6.��1`��h<ۄ)�b�O4Ȅ����b6��3�䙌����@-}&�ݘ<E����{GN2(Q]�����<�4���!�5�;gsv6�z*��F(�/I�K`�c��;��`�6�"��N��3����d�u.nv"D������s��i�K~	���Q�J"g���]cL���Ndm�9�@׵�n�.RhU#�뱲3�CG@� p$xe��=����}M�7��yn{(¯u¯�o6�)�s7rqe1\X)/M���x���������\[�a��(��e5�mv;��X����vQ[[��8f�G
J�S�O���4T�d���|�Dn��B��� �:5�X^5~�S�U�O��{����b?E�����/hRR�8;E��%�|T]�:�7 ��#J���&���xf  �uB9A��Z^�lfSC֌ON��Tą@�[|o�@�;Sm���ڼ�X�k� �����T�Y�RM!lnq�)$O3Ln�'�#ITb���TX�a<P+36þ�21�5͐�h�qu/�U�~/f�����j?��^\�FN�x�������O!<�_\��6J<{[�aj�������B��b9�������*�����D7�>���a�xC���:�q)�Eb�V���T�5;+5��L f�C�l轝���+��8|�)�XALL�)~�N�+b��jT��2>AǠ��kE�ڴ\�«-ټ\�ZՋK��ڤ�w,�>aN��q� �eU̫a�M�ܩ�H���!^p�}C�d�d��֖*�A5�d��_ެ��D�����X�z�9愔UB޺�V
�A`��DqX+�U8������v4#�9&�8���>����Yͺ�;�_P|x��rO�i�C�䔝��H�P���g5�?����{����f}�!��b�6�\�,��U(�
/Y �Q�ȸĎL��y��7�EDS9g����'=��r\���dp����s��l]fh_a��O��?������&�-41��зu	�%�4��n�[{6?l���]�k~|���,��㊶g?�V�28Op���e>M��~\G�[�I�er�\|zd���4bc''�,7`']3������'joq��W>��д�z�'��?�ʆ�t�^�׍��֌S����}��=l���_[E��:�1�a�V��)jc6ߒ�n��vS�]|���K�n���.��H�ZVm��c ��E�u���56�r���~t��O2(�P
�!�I�G���1T�L	��9�BL�_�M�̂� c����_+e�O�E������2}Ǔ�)J1�U���^`�
9	�NkJ)8*>�^����?����?�;i�}O)��� @��ȕ���h�+ѿ�;�S��w=���RǊ*k�J��Cj�5����b��v��mԌ�����Z|'����0=(��#[�E��c .)F�{U�sS�Н��,�Զ������MD�\�#�5�D;�EoY��fBOy�EH����`�.��Z��^��-�l���±C�ؾ��t&�i����<p��\]��j��	U?�}�7�Iq%�>�0�����S������2� rgi��������n���[��b#�g^S���''�:�<���40B��!��㪐Po�"t� �I��l�n`	���uVq!���s�Q}��rMtbPU�,�=a�E��,��&D�d��{t>hNR���^�3��r+�6���%�|{M�Vo�S��"8��J]����Lˢpd�)�T��g�7�n~3�N������ղ�QX&�
���ye����M���I�>���.5	����#l������rT%,�ejC��n��GY�r���P�5��[1A��&j���ZnA�I�ع6���`�̄�ڶ�ǁG�70qV�[���H{P��m� 0�=�@���-3|AA�*����~���-~���4S�����=t��w��F�5��C�?������מ+�2�4T�g˾� �L��-����>��`������MA��>|����@���&�C_�m־��ʸ���ojJ�XB�c��*����������
l$��z�$�}ä鲰1�d��{J������zyaX��8��+vk"^Yjů��qxa�\�gD������X:dx�F��ljr�q	J�p�l7*��V��h(ks�m��\�L���5*��Z�f��-5X!/^�)R:�9s�� <]�Q&q9l��ô�ݹ���܋�R�l�:��s�'�sG���LYz(��8���IpJ�}���D4[�hV����U�ZVź�v�ѮdE��&�d�?��W��W���ٹ���F��~�A��G����eZK>������Q�BE��A��o:a"�^���a2�q����PU�L�fvu�`�s9�{��GI9X"�V5C�²���]��