XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����E8��xj���hm��}[n��P�k]��S2�UP.�쬺{�:%:����|m����H�*	�0��G�A
�1��_�O~������@�0�=x^��8ҷ!��9i�y�_�����Y=Ds\e��t���Y�e ?SL��g�d=ܹ�r�lYI�@-]��A̳��"�8(�:L��XS�m����K�x��!��X3�X�Nv�SR�\y��0_����rM�*K�� �L�p"�����?ph�"�?��jH.�T�~�4��dR���S�<}�3J�*۵��mG������G�E"����l��I3R���=ll����e���50L
j��a�����|��._S3���cn��h}����T��A8���ۃ���!�VSd����L���"Kw�R�XLi?����޸�`xљ$H.w,����#D�A��!���F2�"�[��|M�������cP���� �.�Ywe���~�b_�����͖� �$	�}S�� ��]ݛR��/]~��F��Z>ֹ�W�5FJ�ڣ�/Ɠ�u�ӚӲ��h���z�4���l~Xg��C��>���g�K^�q�M�l��L�`2uR��Hs�NA��7��D
��xJ�q�X9�MVݘ�A�D�^ z�Jg�`i��B!n`�o�U�"� к�T+@b�����\�Q�� ���M2�W�¸U0<⓹,��C�;sv)�X���[�r��8�0,�Q��H�V.*�p/��98U��!�Jb	ҥ�3�XlxVHYEB    1853     810ogF	���ߑ58�כ'�r�.zֆ�mC��_{�ޝG��.�iy����j�*��Dn����Y\�z������~���� ���<Q�EwZ�܄�1�x�b}����n`2�m�<\�#�48�q��A�����\�r1�����֟��%�@�m�G��Ii��A�N�&)T���R���̨���|�.��>2�)��i
��J���3�b�[p�Ԡ�0E�G[3�-�����/O��
�8�$������{p98��'��_�ӓ���G�Ș��-��I^xq}�|�u��3�4R'͍x��JJ��J�"A����i���^�r j7���0=�����d-V�alQAtBa��?��\fr�U�Q��rQ�(��S���x�pL�����듋�-9C̵��:�V~�ndϹ�,B���Bcm���8�9
�
L�`�V�ƙ�8c��cA��.\C��N����#6�0��f��ԗ�r��[1��R������K��aPʗe��@���\a��*��/ BAn&aR�����3ټ=&�i"r�	�hiD��S�q#�%z�@f�>�r�^ݶ��e3��ʒYI�����/�����t>)P�������S�k��sc�c/Mk���h�"�V� �?e#G�q.�^_�^_g������Dh��L���~a�e�666H�}	�\��:��ɲၲ4�����o}��|6�YL�(�������yъ�Q*b�-7ݨ�(�D�F�P�Kf�ܣS��1g�g׻�xCh/5ho��������DW3ʹ�F�5I�k�Y�BP��m�L-S��-e4�(tf�x�5� \ �j�(�0I3C��w*������{�ӼD��׎�>!=������S�����o�`0<Y��u]�5""^V.�*G���*�&��Z�2[�:N�XB0�'�c�j8Q�q��T�M@5?�� �.Y
����~k���]�����
[9�Jw��:Z�\2�����D��Ski�]�ܴ}���	 ��ʄ	�;<^�נ��V�!1�,5c�Т�:��������`��3���ǕV�~\t�����o�r�_kJ��m�\�"}߃�_``=+�Ϻ}�߭\������!R���^G�ტ��n�
��l�fq2&R�/I��Aw� ��jQvxd[��-iK�3�p�@C�_��/Ї0��>� �]�FE��oØ�MH��;m�X�k���l���֝j�
�i�u)���"�WDy�<����E|t2�`��R��w���oe�s)�	�}��ԣX9_���qQ�1kn� ���P�V/꬗:3�挎��������~F�_n^�? E�(0fHtU��R9Ib8,nZ
jE�/.�t��w�2�w�;�W+�`z��wnl�u+�p�<iV�[�����S)�c�#sX�ݕ�H�nR�q�EW��Z�ѿ���v�cI0s�by�};��+�"�68�m���>�7�_�{ρ�"g'=q�
�8r��'`��g�q��k
��]�h6�%f9N��l+�[t��aIg,�ݛz�ݕ��kJPJ�OK�,�+���U������!���\�؅�ʔ=�i)�U4?�u:Ǿ�jx�\:\�&�NP���!i��Q!{�h�&Q`�L?>�t�]k�����×\�S2�REߟ5��{�P˛Z�Yb��e1f�F����	U]!���J(Ja.��2��a�;7{��.4�Gn2W�����<r�V���qIי#�p��I�>�z������8���ղ���dྒྷ�-ρ? 5������8y�<[n������l�AW�:�9_=)�ҥE�B��gn��<�U��v�*@�L�c%�:�x��ss��FX������[��܅�w�i��M��;��<"e�9�������j�Ƞ
�ô���T��H�|%�����|���glj`�21�������� A�������tf���?�l���uq�Μ�I^�5-nX_(��u��):`�ejſ� ���Qn��8���ޓ[ KB�D�I��Go�m��5s�Ǟw�ؠiJ]R�i�� kG��+B