XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����_�Zm��څH�d,��䘵��3(�ԭ�pz�w�W+R��c���"�8�
J�Y�i�9�4�B6�$�C��L��$���sm���?���~��cb�7Z��/�4$��gx�K'�lٝPG��d0d_���H5���](u�6Nл�E���8�⹨�X8�L��������q3!�x�zҪ��tϮ4���#̝�ܯ�D��("���=_͆�-�Of�	-�������o�ZC-��U�'�Kc�)��(AԹ��y�p~�/�(+n}�K�5���� �D{�V6{�e���	�퇵5C3[T�9ؠܞ0�4޿�i���a�5n3�3�QÏԋ���-�BJMIn ���x 8L51Ôkx���[�w�����-�袘,�A�y#�o�Q��z�:�v�:	�:�����QT�w�U�pB�GjTֈ�����v' ��M.ab������}h�oF�h�?�R����OC��ooJ8h�=��]>����B�X�XĢ�@چ�՝�f{`!!$r��'�S��ǁq3�V�	%�5�w	��{��P�q#*�	ï9��s�gGxW&�h�S�CS�A+��-*�/Ө�3	�ґe��O���_�}|�k9d�G���ޱ�3J�u����U���ގ��H�9��L�I����X��gQ�a��X�liB��@x:?��O;lу��tfu�H�}�=.�9�P�F(��;y��[�ڶ>��rb��������̓���[¾�oM�����22㐅���XlxVHYEB    2892     bc0�`,���Bm^H��q��(�*$�3�c���N}<�N��Kv���Mڙ�r��F>��s�3�a5���_ egP
�	d!$�,����TX��8M��H�@bmi�VU�|VO�9���H�a�ن*��F����v����$�J#?�KI�0���v��eR�� �,+*D���WqD<�3H����S��L��A��im��n�6�(�[	��<��R��e��vS�`��k�z��@����a���)�e�g���@�X�p�Z��K�-ӷ���ܥ�ܴ������Q[�]v�M���l�.R8�V�t��c�V2^ô?|�>׾ �y�#m�p�iO.Ll��(	�h���ڢ��U�cΪ����rۉ�w�$^��N%.�	��ˣ�-5|1buA����r��C%��t��7�g���)80~0Ć��5�۽�P���@���q���r�W�X�?�����ƷQn��oU�RI�i�"-aba��?h��m�����v�ԡǲVu�����)K\M�P�P�i��27�?��]yV�-fV���Kz1��R�v8�n���kϵ$���i�Ƴ������.��m�(�4�r�c�
?���jj�xw�9ɠB�~Z�:PĞwu_
�l�2�A���腀ő3��:��������t�H�����.��=��	����W�8�0rr�������7�B�y'�4��R�@�0ҭar1���IhqF���s��&kL��ml��yj%Z��b�+�&��E0� /�>�(�9M3��m������c�x�v�1�:�Dڌ�O���a�Q�G�\ЋO�Շ��uF�D��D�5��T��M���$���Yɫ�:����N���Uy�� ��SC�n-�LX�����~{�O�����݋��E��W�2�����ǑL}е�7�]�C�E�c�GL����M�|�R�,��I�%��S�
G�RO�jDj+H7V�~�C[�o����O1]��&G^m�DN��ʼ|r1i"�_�p�D�}�='q��D
�����u4sa��tL_��X��Rr�
�L�^%he�?�	�雮����V_@��F?�V���l*�P~h���X������29�䄤��Zfpܭ9{�,,k����U�G՟�nd�㿧N8owx9ei�(��i�l���S!���Y�:���R?\�,��Q�����m�`�&�m.ѧʑ����Y������T3}���r�_�Ƿq@�uyy���ۉv�~}���g �^P�%�n�Ǐ�����\���(į|E��r�O�,� ���5�"#���.���G�����y-�Y)�͔��
�:�xyZH�y��W���y6a��9Q{ࡹw�+lC瞻	�|�T �
e�V�82z0
%��ւ��b�e����ء��N�Y�b��E�����e�8TQ����K�2�5����Yanڿ+do06�A�������qB��&��g�o��5!�����H1�xߢ��ǵI�]n��[!t&��?�3��b�#,��%��!Cf������v7�3�E`П���O9��DD���C�)ۡ�9y���S_�I2�dQ�|j5Y4C[x-X}�0��*�ol����ieo��i]�������,D=�� ��H�i�2^ĕ�+n�1w�PT�0�^a#z��ሆ�F�^>eaͩ��	3��)��:i
FRm�"7;W��uw����梊/��8����p9�^�*����hք<Q�)1m�R8��v&��� -��E��W�����V��zD��RDﳟ�1%�m�}��VS��������p�e���d�B��BR�>c|��+_C�y������i@8��2����jk�mӝ� r�,��ݐŌr�0���a㊻#���UG�(�� y�j��k �������$�c�d�KG�l�埰�P}gW��Y��ӋvYj`����b+�FF���^��n;Z�P4�9w��+�*�:�*���������w�vװCWn�/��P\�5v�;���%(ۗö�|:9���=M�l��ä�9�����@7�);t��1�c/�x��%9� l{������-Q�4�S_�ׄ�?�"�@�,��e�_��F�'`�&T�*��|;fbb��gB|=�B{��H��ZR��i0ﱀ���k��K�s��P�ۿ��	��Z�w��ϻr��5�.%����)�Z}�,c���$6�w�K,����Y�kh�R1�j� ��;��9h�g�k���l����4�G����:<�?|���iC\{����ݷ���e+��]��3���%!�T�w��@�����a�|��aC��f�����E���s0>?L���飼zKMoiM(`��&�	3����'Ն1�x�l�^�e��~SsU���̻���w'��9�`L������+���OwUpP%��qʗ��$�ZA��u�����o��@��M��G�ϡ�̇1��#�0;:m<�KO�o�V�����{V�����w1���a�,�/�ya�k��Q��X�Z� N���lߺ4�c3��:��zCG17�Уsت�}��10��Y�"�#�M�70��jk1A	�� *j����y�6�A}2[�5��3
�I�u�����#TZ%�%��{	
�� ���z��$gQ�g9�}�
b�ξ���iSW>���}_i��i|�]O��Dm�u(=!���b�c�%o���L`C/�0��/�	K�>EzX�v��=���� lh�.��T���<�q( ��,�u���3�&��I�9��[X�,��p	��`PZ*$B�Ψ$�#����I]��`y�*U;r�B*g�3�L*�'��=�RᔖN��r~�O�d%�_pQ!��	.&�t����G,����x/�&]��>J�ǀ����ɟ�O�a��ə�8b^5L���e�y�}y	�L x��]�r$�h�t�BG�墸O��_�(e������/�@"
Z8�B�