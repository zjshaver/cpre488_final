XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��A�X��&�R�/��7�)�/�	sJaA	<Q"I��%A��m�u��6��S.ޟ���O_��M��&��aw���x���NЃ��[���A�H=�$Q�<�ᒞ�@�z����$g޷�\u��QlⷠV��MǾ4��$�e/��BĶ������☞g�?��ߐh�w�(]��P</:����+�ݞJ�*���A^D�.9�Rx��P=+���+Y�	\r׿!axB�o+�EQÜt�����5r��d���gr*�7��gL�W�1�^x������Z�,�/�l� 2OW}A��X9�3k������������Ka�[�j�����pF�3S4ۓUe����2<��SS%f��+��ь��G"�u�+�!���J�N��{�W�|�8�=.-��Kʑd͈;�PU�/+�Ch&c�X��̶�ܢ��0m�k=�^���W�����"�*)�����4��͟�¯1kx7(H5o�G����~����h��ױ+��svu��kkL��ؽW~K��b��o�ʌ��sG>X��&���]��Ȝ�U}P\���p߃q�ƍPl
��p����VO����>�T���T�n�^UKw��P��uϺ^'8CS��.��(� �>3���-�dz#�?5�J2��۔�7C�`B������Q�p�C�i�_0��8I��^�� �m"��C�;"�R~<#��N*�-�@ڠs턵��A�<����G��L��Uԋ���	)f&�2� h�ɸʊ��ɘ�A��G<� Q�XlxVHYEB    4b9c    1300Y�����9	�4�#�_�����7��y lf�i���,����It���� �������"s���-���	��5S��ZL"j��*��je"
	*T�c�7�&�5(�O�JT�����A��9�sn?C`��E����,y�ț�f��֫�d��@I���T�(�$s�nmEU�n;Py����C�q0�"��C��!��A�1�GN<B�$�Q���n��/�b�Q�c=[����£��yop�5PDg��P6��tc�m;���%U_����:H�<]���$6�#j���jK���^�]�1����=��P��Nr�-��~	�tZ�|�}.n�.��j8�a)����<�0Dp�@�㣡K�"[tw �pؓ�����M�@1��K��
�]�E�OKq����ľ���3���:����,]�-2z�*�]݂/<5u�G~�D�,����\1����͙�is[Q \h�L�eB0��=�e*q�f�GJ��ly��3
QsÇ�x����m��AP"y�]�5F�@�A7p
yʻ�jS�jg:e�D���,�����0\���K�PS�������*@xi��^w�}��?�W����j�E�P�|�ƻ�K�������ǐ��T��0���q��ښ(����{d��3�/������ZSsړm���M��lU}?upzP����'$t�:|������=}��{�Ѐ�/]%v� �#fJ���s�������������Z\�!֯������"��}�i����M���}	>���aX�B��� �퇁����V��e���n���I����uY��C�[�ڋ����\� ѫ;>c��S��P<��A϶3��w�D��}��'S�Ki|�E%a�E�)|�������5��tS�0�� �Su���8ƱMW��:�R=��@M��Hj!lyJG�+G�?����E��Z38�������Vu��oD@@T*��
O��{b�:^��<�]\�"�oVez�y_#�'Yd�%�#��� ��\�����%�K&�ƫc�<�1a���g�߀���i}F���t���nZ��I�5y&�n߅&`��
W�W��˙�谶��l���*��2�7'�K�����I��T��T0�ltZ|��dm���E;sH�`.�N\i+���G��L=��=����p�gƟrBm��Z����L�h��G���0��'�>��`F�B�C�k�!E�=��#����U��Z6�!n2�Gg公��}�rn�^)���^�x|*v�C���7�Zླྀ�-��nĦ��R�)��o.w/槖)�Q��<����z����V�.��[Q�22{��]2������l]T:�6P,���5���O�B��G ��[s�[m�6��<�ǵNԪ�s�d#O�n2,�3�͒��ӯN�����4�a*=�ޕ��'`������9��.�%or�*�7F*f+�t�n���e��B�8���#6�4��e��X��3:@tT�+����b6�9�#��--CT�ʋ���`�&�_0 t*�!i ����5Α��΃�G�r����H�7L��H���3e�%���4�޻��T�do3�����Oae���k'���4����L���ȭw�
-�~�G�dĲt
��ƌ����[�̢�T�yM��c(���"J6���=c�=�]�H�T�Nu�I��Q}E��Ч1k�=��X�u����r��֜��,��\F������t�����d.��B�LD"�I�IVL�d��%l�!l�[*�Uo���=��s6����eFPdoZ�ϊ�a�r��W�A�����U���j��r���P�k���j"\撬E�=&1�+��+�TP�h{{��b$R$�~^n%�L�&���3�}�1�۳����Omܑ�4�^m���J��a�R>�Ƴ�q�._=�O��r�{����E6� ��O������4B�u����╧?�y�L$hAn���0%�4f�6�ز�w�'���8���~K 7X[c���~����r�ū�uN�����e�N�\�w_~,��UG������閱#wyFs���W���/���Iʮ�����EX.��O�6�8�r"��w�te!Y9O�~r~��_�aS���=�hX4�P'�
X��]�ݮ�����#��5r�W c��&��i�P��A����V���n�Xx��"��6�s��"�7Vg�=����&~6ey��AP_5�S��5���G���䆗^5��ϡg�b�ٷ�9ݗ����РDńYFJm�0(X"��.�'2���XP*3֦m�t٥�Hg���#G]fj�KoE�[���HH?o�����˩U��� ڲ�!��mا�'���nWv b��r�yiz���]4n��2�g}ð��	��66p@S�3�i�ݕ�M�Qd�XV��6����6������$�-/�V�)�s�Խ(ۙL�Վ~���JHx�_���u�gϽ���;!�A����]�=�4�)~���ڂJjׄ�b+wg-�Cx�哘~�ǏW ����%̫A���xJ��qr��翄Aw̖$�g,?��a��0N9=z����W��ې�L��:Z/���#�LvB5̩r���{���|!����[��<S ؠ�;3�*����ū���c���0�����3-	����%�+�?�OR��c��C��-Z�'���ao%��pM���p+��Oy���#ʚ��>uI8y��ʕAr�o�ig�ua2�����F{��x�bx�SX�H��(���]��$9���
| h��w�*F�I�ѫ��0�ܡ����E�Ӛ8ŋ�C�N�.N�\H&����&J�%�1��ڌ5��֘p������&@Br.��Mu2Т)�F�4aI�{}sk$CUw�k�3�z�ys
�C�K�O���d�`ƒ �0}Z8��g5O�&fU��t�AE�u�������?�*�{�^E�G�8����v�6	sc?(�m�7�F�?� �P��?���j#Ǎ�?�^j�l�U�ƈ��C���c�N��&�Q:Pa��$��;}�S���������n�� 6��Ņ�$y��Q�<�ؙ���Hr	���,�ʲ����9��n�yl=J���<�����,z'��2W$��ү�U���	�7�ȟ|�lڪ0�v]�f�G'�]���⤼⚿Ӎߵw�m��+L4ph�J��$Y�0�iJ>)�!#�b�~���Z�`�!�����>+��<�����o�R��P޹������X���v�8�nO�y���|��ܙ��Kz�=}�X�Q̻vbn�ߤ��V�?4��Ϻv����֤���x�9?b%6�{�����2M�T�{�x�����\,O�� �hLوq�(���:�f��t�s߇��;�߽CN��/B�?�3�s5F�~c�D&P/B+,gq��<��f��\�;�E'M���k���P#��D�����z�8��ҡ��C�V�I�NY)�PҶ�&*�����-p1�d��G%!r��HV�������	Nҧ �%�ߜ�i·;��gK	���Ư���t����-�F���=����=;1Eb�i����>��P&��;-{g�������m�$4���B/����b#�=���������Yi�R������ߤ�7>QW jp'@<�� �;�b�zrD�����
;�6�p����"�
�sX8��2h;�-Cʢ<e��$U  �.�rq� s� ����#��TtN�_�[�UO�媅��y��W�L�cy��n0ܭ�+��C�G8�F�u����H�bMi�A>����af���̓L�TJ ���"B�kb���]���<��@V�#�:���� =�q���,�����ӎs�p���}-����Zǟ�}
8�+!��I�M�:pb�2�`�6s��%췦��*�
_$��b�M��ɹ>�����n����L�ە���8�F~~�a������.�]�L��O1U3�����H.��Z�>u����|@�i��6�q�cP��
\��ϲ*h�-��Y=ݫ4�CY���քS��������LHF�&�$5��ze�\Z�./=<n<���E�iШ�9�W��,�9�'�����nd�Lm���Lm�b3O�tH�{�'�T.Bn��S�� a3K2� ��sN���kLT�cG�#K�x��ƺp��MpM叚t���{qhh`�O!M57�H�="Q���ڢ$v=�2Lb&�_(k<+=�y���=6�Փ���,��_�Z���"��ӥ�m`lX���
%_��m�v��`��6vT�՟�R+�(n曄������r��a���㙣�ƽ�����@��FQ�e�2�=�K�"�i}�1��R�7&�����+{�c�|\������H���_�ϿJ�_��Yd�����#F��Ϭa��T`�BT�b/�����n8�s#�����/[(�Ӌ>��������[4D'����2���:�(?{GC詚�hϻ��<�37G�f;�d��J޲4� ���y���9OYZ���S)9ҫ��L�#b$�~S�͚P���ܡ��!�u�y��x�Oe?9��NH�uh{�nn
/L��a%��@|A�/[��x����*�����(�=�M.��H�)�H�5�עnT���ǟc�w60��~�EwQ>J��n���[i	����j$��b4�{&T�'z�s�r��/V@e~O�kFFRT����01��]~|�%3����O��"b�4j�sg{�q��L�;�o��/5��I���i�4e@M�2