XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��X��x������f�ʑތc΁EZ�+b���]�,ل|�
���F�Q(_;S6m�W8�'a�l�.͠�G��$�s�fq��$�i���@ͮ��>,L'��-��.U`��,��ܥ������ܻ(���"@�~H��}:a�ۅ��Y�u_B-�F�˵�)���f@=������NLJ�(�B�2�I�}hEh���7�|V��j<�LӘ>Ei�{j��ۺ���s3��� ��x|sQ�UB��+Ε4:�+��������T7���{�aA��Md8'��n����U2��`e���~n�,���ʮ��r���$pk�ݤZz�������G��tZ!��QG���N^u.��Y����/l�����e:�
�����U2�5�7�k��V�Ӆ�=�B}P@\U"�P,u9�m?e��r}$~!/��~�/G�r��0� N.	q[�+<T��d:Cn��~,�Y����W��j��c�*!A�T��j�	�у�3{ ��^5;e?�51��o�`QA����ݶH��\@}/9D�n���8�d!.����� a�!"�!~�>�M���.�.{[�kmLx14�]�\&T��Җ��w����9�^�m���~�<Ŋh�k���,��K���D��{[��o��cp�9�x�0}#�O݀ljϨ�na�$GX`�.x�F�NR�Ū_p�3����wF%ȓO�3���
v�OZ�(��:(���\��96d����i,� _��o2��ee��׳	🡾�Q�}5�_F�O*�XlxVHYEB    2892     bc0�=�	�Z�S�H�{޻����}��>?�B�Q#���Qog?�DNH�qý&�*��fװ��� ���R[�{а+Z C�6��j�%�p���8�8T�x�v��+�)���
l�뷺5Q�1��ύ	� �χ�:nIw��n�_H��2/-��s+�U���`�d�m�#��r#	�������_�~���S CEn�0��ʗŕ)=��RVP���%7D�Dp'��������/�{!����]�T����㕞4:�%%bGA]A8��:~V�����`0�m$���+�:�0����Tˀ��O8d=�#��&���Ѹ7�5��B~~������+�5�.���t2�cq,�;��9��"�_ߌ��z_�=�:�����u���c�e0����:�ƭ�(t�%g��b�q���g��.�W��R������n�q�C��!fp:`s��B��88�I�2��$LjU=�����Z�e�ݱ2�jG�4�G�fD���Q�'M���!Ӽ@8z��>��A�l���z�7��=軆��%�('��h��@b?jU��������ƽ��8����\,G_|6<�P���~�UޒF�J���wI
�|5㉆d�(����0�`����ux_��|������;H��ս8*7A��zM]���D:�f\�l��b����[�"��ՎSDj�ZD��4R�/�Y֭��0��f�4G�[�YP���/3�����0T�ȯ���<��0�����&y�ٞ��?I�349/.�J��ś]���;���JC�����h����'�0a��r���5��񛢊�y�D}�	�gj,z�DA�Si�!-�o@ߋ��u�"Iӂ�m������ ћ^�e02ٔ��%2@��FM��R�8'��$�,��m+%��-�<w?Ƞ��Z3Z�� ��*��Q+}���z�� �Q	y���;�'č�r÷5�q�)�}��N��P�k�ҟ�˪��K�o�
�� �[8�恹Dݡ�Em��M������� ��ׅ���[��)w"����TL�8.ɱ�7'���:�P[���=m-��]�w�5���K��� 
t�֬�L�C�b}�Ջq!5��P)0�}�@����̉_�7�c/��MEC��i�E��8��K����3%z�i6�hQ���{.,������Q����f��JH<n��� ��;���>��l��~E:W�l����f�Pf�8�}g3g�+h-��Q���5�x�ء��y�?�0n��	�%@�(��EQ�� ��7�-�/W�����S/�d1Ν'��S�?��c�.
�Ĉ��R�M��]|��N�!��3k�;��=C�ZM�/=M���B4�R^R���K�e7c`#@����<4��;o��m�ёժ�JJ -���
��4�!wxi��j�����[VF_ϫ�2�Jn-������J-�[>#h�;%�9V��&ݣ�څ�W�u%��jvK��,�$�DRGG�s���N'z�g'���E�k�A��/����k_��fj�m'�.R7G�T��ɇ��;�[�u�7��(H"ڃ8Xyi.��h����J�Y^�Jc�z��l�gӒN�G�]����՗��E}��PB�2�	�"FR%�� ��d��9׾!qK��+IXp)�sf�M���}A��񫐂��h���k��P9���X��́��>DI����̡�og��z`�߰٠v�k᥀��њG�v0ï*���et�|���HFy���}Q!�4>��S�!4��w��~��Q�d��������>�~��}���:Խ��<�L_z�%1\����⚚J�?�߇�BL�Pp�h���5���5(B!��S� ������v��z����O��V�\�y�Q�o��vܮ�	/�X#�mI�zd�����W����Qę����Hْ=3��l�oҕT]�� ��B������lT��.�}���-'����4sb���;���Р���03�V��������B�m�`�3�& t�ΐnW�nr��"�{7�W����^�,�]
t���7�Z�4ޚH���d%���5d���|3���+�*� o��E��ie1�Q�8E��9]�%$t	�0X~R�R�Z�Y�	`�����PP�I�4�y��Z�O�u�b7����,[%��)2:��"���+"I�����p�Ttz�d7Ly�7��h�@?�M�OcAP�i�MN�7��Qr!q� �v�`�q�3nlh ��d�n_�
O����X}�|������ ���\`xy➗�SU?�&�}dx�C6ƛ\�A�:�1�i��0�dAgY:��{��pRxБa-�*w�E�1H�Q��%�M5�>�����5���}A��m+R&]����N'ㅣJ��h��!fbQQ��j�)��E�nt��%w�=kd�*�Cz���Ed쪒p�l ���p�����%������rd��$����8B*~������2
�_��7[�Y��T6�V:N���Urʳ�)$��HU�ׅ���֥m�[��u�Kߦ�W��R���n�jm�yu}o���T�v����S�]���*�T��d&����t���o0�0�(mmP�8Ib����;'�����.������Q��?OF'�M��]}��$�w�5��"^Ve]�V�ڙ���j=��c^�#���y��-q�V�~Hģ���M�c�p��=��c�;Y�s����;V��vrn�����/��P4��8�%c92�x]�n�cAØ��/��(NO�H�)� ����t88�*��a��a1ob�>��ucE]H~;�͉+�d�F�Ц��_��3�M���[�}��S��Nŀc^�l�p��+��kY�c��˩��	V���S���X���A����)���P��ݰ�=J���t�k��;¯�����5���Y4- �db��f���HdL�V�����������:#DhV����d