XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��x6)�ܷ����m��j=�O�h����JcO�&���8�.j�����n?���Nҙl%�����4Ej=�~����tbs\�#���ǎ =�qf�}����"f e����+z+S�=��f8.~�0!R�fp%danK���^v�I��������-o��¥������z����I:Wl#�ܐ���tKxl��M	<9{,ǁ#wbci��B���c�Z<� ,|m#��%�L ��Md�Y�ջ̂����K1����� e���$w�4HՃ�/<��r,?SO�9��`Zce��$%>4��[�O�Ȣ  vb���T���?�NY���P�0���*�-����uˆ���i�� ���2 �>u:M�BV�o��M�J�GÕ�s{yg�ma��6_�2O����67����!��d��r�Fݱ��{x����^W��F�0/�����Ԍ��w�$�dX�̝�̿�@q�5��ט�W������;���Q�uGK?���Ǚ���N�*p�8������{|��"��O���!��V��3Ϗ	�$ltv��%%>A�.t��Fy�z�1G�.)Nqbת�ι�DL&.>�f�hKL�%����4Ȅ�zN�ݠ��m�eğ��p�uw���*���j�*Vq�7ZN|R<{E��-�'�թ�����h�V�^CU��c�{�k�M����.��4T�ؽ��@�9�๒Β9Z�y��oS<�m�,���v��@(黿A�2XlxVHYEB    17d8     890���J-.�c7Z��9,β+�x��,D������:��^1kp�k�w�5�n)�u�i� ��ad*�}�j�-¦YJ
�� G�7q�"(���l�6	�B�u�iqG%��i�5��{��z?�D���N:`��cQz��w�W:�,8��eg�B䯮v]�N���Y��O���6C�4&$PH�;G�5ܱ�)�z�	7�|V�b-������w)�y�[�d�2<��h =�oH��N]F׉:}.����y��Q3��Qb둘&r�v&qf���ċ	_a格OPh�?�&0И]9ǉ���p�6��S��hB+}|@R ����݀��yu�Ƒ�k��\@V��Z��ڦ)��0Up!o'~�����)g f�tu=���r6@������e�D���CI�׳�^�����՜�K�����x1�Z��VEA��̬����c�8����"'��F��g��?h���;��̭
���S�Uơi@����6YŬ�$x�����ښ���ɩB�=��awUDw�t�����o�h����PJc����k��Hy�D������`���ǏS>e�!P�tw�G�p�F
a}��w!��s2f�6�=�Pz��B�.G��v���[����0�iQ!5F4��@SXB��5�N3���_��S����3v��� ����V��{Qr��;��,D#nl�o�++�.�n���}���o^z�Xɐ������Y�V�bD�U ����A]an �GA>`}<��_�e��d/]J�[�|(��������{�#�п�@��I��n����L�[�j���I��Xҁ��]��Or�d����%"]��c|���	�8����LW1�u�����ʥa�wR��Dl�R.n�Y�\���N?�8��:K�r�֙F�2z�i��ڗ�̊����n����.%a2�҆2dԕ����X��x�m^\3R�c˂N��+_�<p���:x��z׊Z�;	zL���_��n��h�Q�pv�Ll�0< �r�X[7��/�==Ku����t9���Kl��?�d�,{�g&wl�b'U�!�e�J���V�&Q�~n ��v��
�_̌�] ~
�i���O���Y���5�'��
S;'���'�>iy��sc��2K����~�2�X���3
�h��}4�e��/�f�ٯ�N��ߋ���'7Փ��*�e��<I�ȿ'�E �@ORe<�eb�ú�}�*M^K��Q��T/��Q����h�|Vs�_��ۍ��j�"�/!� @F%����^��خqGY 㔆�b�n���m5�Y�����v��w� ��g����k��7�K|��7�e�,�n!Tbf��a�7�\ш"!�"UZg��J�v:�����"���b���B�� q��r?-�������S��>�k�rG�`��5.l�����8�JP?��[\�q���'��hYiF�;Uꬎ}����@-_����\�v-��s�	ٺ�:$m�Z@���&5�BT�ѣ�*�a��kD k�sni��� �8����M^L�y8���]s��͵=.�ӑ/1�`d["�J+3lE�O��y�6!g��T�c��Y��/�d��ˊ����(��ȶż���Ԭ��[��if1�}W�$U9N��<6���2��!5oӞ��E���j�pÕ��t#c3@��:�23_�5�h�-���2w�~��晕��"����
O&⇹Xu��;6��+���\zG��).��+���m��}DZ����M^H�n�d/ �H^�TPT�?Xޙ,�(�
�Hq).ɋʓ��@L�nѶ��K" �Y�����>��?�K�4��M	�f�$��~�_��E��\8��8W �~��9E�R?B+s��'� �'s0J����jP��V2�M١���vV�a�B-g�wj,e�1��MVokjȆ%	=���6�{��,��[3i�s�'Ch�g0� <��M�+N�`��jG��39?��v�)Gl�f_h���~��s�|�ğ�����!�ڐX��c�B�v���I�toVt��FFr��(�io+!܂�kG���N��ZO�D��{S�fO� D�� Q����p�~�
w&��cU��Fry�Gg����,Fl��,}�1����b��1*
�wءD���V�^��