XlxV64EB    1c03     980�Uݑ3k23FG��@�KE����[t}2e��"uRoG��,����a��՝ϟ�(�7UJ���Lo����7��%C��9w����5Q6��<���G/$\:�$s�;J����X���| ����Hx��k�2�uaƅDRg�AO�)j�+�����~\�N:�L�����3�IB�Z�7��)���]AGy]������u���孮c���pb�O8c �@M�ܠ�Y8�h�<o|/m&�jD� #(-e�p��`�Z|F�P~�0�
���u�XB@��2�������ϐ�h�mv���DwD�u������b���}�0���Z�KLJP��3�����r��P��q�Շg��p:m����f�n��A�n�Zc�t�^��մq���3[/��o<Ͱh�r���l�O�`=�&�يT(�hMN����X�e�?�6��ER�^HP�x<�~"�2#��&ǂ���ΜT��.�r4����Bap����㭕����X�����t��T$d��m��GS6 �?��|2�J3k��l"��B�U5����zf�WU�퐴Ş+\���;��a���~;6��^��䡩���2j=K�G��(��@3��/�/3����r�x��8�3�Ý�����1(���ҌϪI���W`_2�:GP tVӜ>c݋�}8g�����N�`W*�V����%�y5�*��\���t�F۸���8T>�1.�{��%w7�@Y��� ������Ϭ«��ϣw_��!�����/����x���ȋ�XS�u[s��N� �3z5ε\��3#}�5-g�h !ֹ�z�1�6σ��^�69�A�Ay3�� s�/���i��"p�p�!����{�O���:[%�FDx�^%�e�,x2Xw��~w�;w?�|x^�b'�~]`Y�<�h4� 9�:���r��^�������~G�jw�`E��J���E���k�1c�a�Va�\ �3\c�#3��ObA�0y5x�p�@n:>������-���b��AB}'��a�u�eV��><�{6����Կ�ȏ�6KZ�7�tP5w���֕�\K��<O�SF3z�?Z&1��-64%�a������~�d�٨�Lb�K��-^Y�PA�f"�
@���a=���5�4ԗ������G�4����L9	��E���Z�mF��]"f����X=:�S.P(=�m��v�
X� iI^�������v�#�Ya��o��-a��j��M�w'f]�5A��+�ž�IQ\�D����VJǯi�FG�{���hO���ӤHj�zT�;�`�ή5�!���P��+X�8N`C�+)_�C�v�ZǼ�t(��L,�22��A�Tz�=�\J}�)��R/�dE
�`�ہ��A'�1��S�a;�Ji�غX�-���l���K���	�ؚ�/�N�:�u*G��� &��yc���Gwt+M������3�Z`H�I�8�mc�.�o�+~'�J�3!0ER���6�nd���ߖ_�O�J �K<� �u�ס�;�R��M�'aﭳ����K�y���`�/wo�7ד�t��}��j\pc�8}`�g����Fw�
��	��U��	_�W��Y��j�Iٷ��N;�� ��am���%2[崸�ogG���d<[P�u��Ol=�6�Y���w`����HD�s�J9&�%E�(�-����y�A��*�l�1���W�&hUk�~ň 0��W���HT:�:�V4�?��A����)��Ǣ����H�E��wgQ�#��A�D轭nR��r��y)�/��d�b�������
��=���!��I��9��*�~(q�ѵ��E�V��li��?�{��C�%-��w�为aed^t���赭��F]�t�+�����Mn�8J	��l�����'�����k���%�҇���~F.��k��0����zҐRe�+rΓ�:s���q%�]46�R�4"x����AV�����1a��;��\Gӽ�t�ԟ�S2��A�"/��-�����4}1�(�?�MAZ��G^u�˩�|�!����f>�Z�G��,eŵG��Fw�;���tyU���$��l�:<���〈pй�&2���ʖJN�X��������]�E��
8q]���j�㡷82-9};*��*��˧uujP�j�J��$m� bX�O4�[���6�m���M?�u��al�sN^M<$P� )8��S�Q,r:à.
3�-�_/��	]����Y��3l�6���T)�,J=/�[�ƙ���I��C 7�� ��lt ��c֖m�'),��W�!x���.�aٽ��du�����_lΙ�gkB��G��Cv�ط�*+m��X�>;V