XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��V�y��Jt�O�΀"�{P���4�� � ��f���&kv�_g4/�l  �81�����Q���[.m��5�lw5jd>�w�|ׯ�}�_10#���'W�h$�ȉ�ڔLBz.+[Kjj�o��D��uX#����̃���g[AԵ�WYa]nh3^��[hN��^����A�!�l���=i���F*�QB�U1-� :F�o�R�c��s|�=�M�S����u��r���[uu���y��译S��	����C$����Ȋ��pz�lxo�(��-�Z�� �:���SC�ʹ������	���W|��k> �h<x�o@��r)�dV�;�J�qo4;^O�IENٝ��h|�I���p��h�hF���lC��QD5�s��i���p�}Nu�I��>>��ShC��$�^���'[6[J�ZUt6,���� n�P[�y��V�A��9U�r�� )'��
�Q
�ҹ��v`,���S�I��Es�f����2�^�x=�>H%�9Sm�1���[2A��s�:P���A̿%���R��^Փfd%o?��\��kBq��4L����s'/�w�:uQ�@;��[�\l2{_a+�M?�Pv�er(Zg$u��n��,Cres-RD4�3��͡�t�3�,��:
7&1��m����r��j���:�OWY����Q0
R4��&e�tTo"�j�GR�?-�_(���H��hd���x\`}^|I���C����H�m*�EI�l4�XlxVHYEB    70a6     b90��An��;�ѽiS.51횁���(����b�e��{���ǡ���m=~��	:����n#�!?�y�/9Ӫ��6oA��I x��^�=�T�3X�+�$�uk�c�7����u�}��4��'�]�=m�\���	=[�1q����]��r�8 a�Zv����(�)��p�d8�M�M:p_��w��9�t�rWҦ��"�ԅ�07���>6�m �e�HG��ߓ?*|�5���Rs��yܓq|{�B6�J��"�Y?\T�&���+����k'4�>j`C�/�fK��D�����=`���joX�����?Gv�ϸA��!������c�l���p%E�z�KoNO�-�6�N����։9p喿f}�����~'5���+$�`��0\�"���tBKE~Qi?5�� �)��ӹ��8�댏NѬȢ�Z��n6���TL ���])IpMR�r�"*�XU3�q?D�7'�f�Ν�X�i�)����wq�]#ɕ��F�F
au���P���Yp���V+|5�%������ ��2	N�|{E^#	_-[�ۿ�7�U��}_��ju��wy��6�y��x�
s���G_?�����'�O�'�P\5����C����T|+�XG+�8�M�}��W��G�Dr�,Q��}���7֞�]p�R7�.�L��r�?ļxA��u2�侂lP�HBZ�'������8�y�`v��Q�E���5�<���J]xWyD�\L�=�ښ�S��T̻4�R�P�./�c�5��i-�(���%��0/W5��-�� &V��Q4}�,9�9X;�ɵ�,�q��#�o>��*�B���ы6�L�~�����-�5�R���*<�]�����p�L�*�7�#��y%����J״�䎗����Ā'�8=:��ܢ��ꭴ�Qd�ڹ�����V��QM��D�9ɺ�K�C���ź�p��͐��$�`Y�BP���l��_��Rsbz����R~���Ͳ2̋|��l��]$4�M7��(ƌ�3�˺�]�Qv�YQjR9u?�uQ껁���_������.��Y�s���t��L�H��T� ���X��V�Jl�j+�f'�2����.�S+a�}���S��f!X�QW ����#ϐ<cw��s*,�S��I�P��"�������'&��]��cz[�C~�#�� ��.��l��Q`��v`�X�	Ke,|o�NZ��L���A�Y~e�d<�sxv
��K�A�M��"�"FA)-m�s�<w����N�P#���	��Bk>cח9-\w>a���=�w�^U�48 T�Pt- ��1q�Ir�ى���NW�y���|��^P��/�ި�J������͡�0��¡oQ�|Ǖz��̐W5�|4�w.o	����ԢY�w�S�?TEǴ��vJ!���#g<4��Y5| 5��ub2�ܾ�@(�L��Ho��f��*6����>�-��	b��FU�͗i��������_�{;<Ff�@��<�����_EL,�>�I6�zM7o_ �i]�;��E���/�|�T���}��>�A�Z��j��&�h��[�Uᯣ 0��\���W�D��t����ر�}����~�*�zs"�V��p]g�?��V�Uj8�J��R>��W��i��8!OG�4Ks��H`�+Eқq�l���7���u!:e��L���z�UJ-i����E�@�`�&����&Ֆ7��9)UF�G� ��Sp}��P�gO��f!�U�	n�i��S�g��a���ـ�tݮ��
�F6�BH�?�od�K.?�7Z����[DY��h��@��ؗ�e~Ŵ12���S� �E�R�6QlI9�Jv������7�[(9s{����R�Ѧ\��۳�|�(�߿U����װ��[Rr�,je��Q� �c�<Fw[�����������X�R
&'��f���cR.�kX[�,��f����R��4������='~U�%8�`��8��/����щ�JqAI���Uh!��N*xc����um��_����!�*�C���-�jQ����_���x�2��@gBa�Y�8I�p��WL+��Us��f����$4Vn����/�;���
�^iXk池Z�aϢ���VhE������{û��cg��Ut&ܬ����t�b�~���u�s�P��*�%�� M����<ܒw���������q��j�:�Ŕ�r��HP�=g��x��\���=<{�������D,��/���T_��ng�z�����\sS�g�9H�z���B~�q�5�,0�/� �U�)i�q�a�@?��2/n2N�9���ޠ�Х^[�DC��c�f�y���wz�r�� �8�-�G�D�m�,J����؇� �7zr���h��^*i .#ْ�\M~͂�ƟQ��<Bg&�T�5�m�4_�̍p����MY���$Ȏ�57�*P�iKB'���xb'�ZId�&�$(�7��nGB	��s�"�ʌ$�L��$��D�A))�M�P�~�^�?-*�=�� X�U�{)�5~&Ȥ3�x�-�K�i��*�(��U��C�Y��g�������И��h��|V��lT+|MK�����2��}۸cr���E�Ay�5e`)���%Oμ��^��!Sv1@��߾���W���	��� ������F82{�4%#a��@����v�WVC!׆.�)aE�Sr���gF�AS��9��D�ű�C;��!�y�ww��*�/#��dw�����9��l��N���JX>8��٦�ɭ�(�u#-�I<�/U��!���7+4���_xꄇZ4'צ������l��i��eT�c�`uy=.�ό���R��%y��RE�u�ͪ�aD|:
�sy\�p]aJ��	ԝ�J|$X��;��8fjk/,Wb|:��