XlxV64EB    3fdb    1160�-V)c9�jN�t�&
��6ւ�D��5��o�ͦ�R_�A��q�0�M�y�@!�V(�8<Y��I9����;בCC��&��:��ȉ�w���8Ȳ���.dB�@w"��O�� LQ��;��_���\�MV}��P{��L����y�kt2�f��%rXw��	<1 ��\:$�5�~]TF��V�NSJ`"��,ቘ�����k��$�OG������ज़\���M�0ls��S��rǓ\�����dK�M&��]�<|��8����V��R�B\�!Q$�2ֵ5��;���HK�=��"��("f-���
P��Kކ{aA	����7�����X�X7���p��Rk�G;�ǽ�C�����sX�\mdO�8��I��e��w\���ll����%�s\�H^��[�q����3�_���?E0/!�X�v�ŵ��˓ˤ~on�v8&S�u7�u�7ֵj����&f���n�<�x� ����E:"	�G]&.s+>L����>r�=k|IgEk.�����:z7*jc��P��/7�� ְ/E�1�c��X�����9I��,6'��bW����e.��%��:��6�G�p����D��!�R�WǙ
��&[#L�)V���*�|c��F��1V[蜪��?�D�@UA�M퀴n��EiQ_fG�K��0Bl8�UE̃�q�9��/���#�_��>�X;$z�Ý��mS��U��D$�e�����zwv��ES��U1�*� Yb���}�s�I7���32�� Н�9��}L��W>�����(Ey�<0��$��bu5�>_ֱlv|Pz-;�8j�|���QVh��Y�l��`�����,$���ز���j ��K��n���,O��(�umX?>cE7W��-q����>&@V布��?� ?�M	��$��#����费s;��+]o�u۾��\*�j�`J3�M��h��h^����u�9ĝ��ê�xdn�P�p�8�@�]�U\k���9���B<�����hp�$��˿Y��8)�����:��2�WV]?���إ�<��>d�F��K�i@��WG�71|�,$"��=�X����!�X�� t{�����g�)��b�7��Y��;R>,=���-�7_��ݒh�i��&��Px����b��P����S���aA��_���*�5yC:�z��I7����t��A[�X�ԑ�e����b<,>�]!�XߕJA�����ċg��/X{>�K����Ε���`�	�r�Lq($tJ~\-vK���g�n��U��e�$��SwI ��]�Ɇs᱒KBl>�<%�Tn~���l��R�g/&�y�lӫ���j�R���������SO;����.�G^�0�x~�J��e߿��V+V���Gw�Ji�������&g��L��k�HL߻�ڜWh �x-\��\��SO����	�1�ҺJ���f��KAR�>�.���te����Bw��D�#=����a[�V���~�
į�ЉI�M.�m�ln�1"c돻am������̥%��~Q��!�b�u�y���ymdN�#���Lz�&���d���p���Uͼ�D)�[?�/��K�,8��2���#fȀs@�lK1>�����u�=�_6�S�3x��RI�P-��YƳI��?9�X�3�����X�tɑ�o���:,��' 6�ǈ�e<�m�������ܵ���\���0M�*�6b���
e�I	���.+1�7Z~��[a�h�gΪV��c?���b�0�Q�=\d�h s�)�)�Ӈ'8kM��J���.)L'�F��"4lƫ�8�1��K6�<۲.�s��ь��s�f;G/x�[Օ%�ˡf"����5������3���0��T!>�C�F�Z�ZP����G%�65`�d���A)Z�
	r|�Aq*Z-ɣ����_e�� }1d�2Y�깐9K�����O~�k^��j=��_�z��r�2g�~}2��;[���O��U0<�ڌ�~D1
c��y~��Y$�qmd΢k� �t�'�H�u��C��5�� R��|E��j-�A�?�����:q��˜ß5 k@1�o��s��7��LW�N�0��#j�h�T��R�����|�Cg�ng�?md`���3 tI�d�D�Cu�c�-�1uhXӖ�.{���y�"��f��F�O}� ���h6�񕴽��_D~��]�ao��#�?�Nd�h����o��y��L�C�lJ6�PeF�p��c1_�3����jK�-������?��vbѥ��tnJ�(��o+o��?\ʋe�	r�-D�ܵ)p__+6���u~�*��	�G�1��;y'�(Z$#Ҽ�>j�����OFxibJ�rN]�sߖc%�����\¤�Y~��8�|�HE����v�����X�8�y��~�?u���W[	�2v��7����ܒ.@�a��qD�>�hX0EER�ͤ�+�+6P�0�S�p��c}�ACM�y^pg������ꟕE��+��T|�w�:nա����[>��t1�8��"����k,t*'H��\�nC:����i������)��V�}�G�|Kv�7{�N�D�kj�Vl� v�/!TK�w�h��A�,f�2��g���֖���[�s���W�)osլ��rK�zg����rj�tpd�+�@��Z����̧ؿDH��e!��5���9>џ";HٶWvb�����R� 3��Լ�h�+5[<�q���#��>R�ɟ;�9o�̩�ݫM��tb�>$32OR��ԷR	��G��ܵ ��Uͷ������B��X�z����l0�d;���ol1)�x-�blW��� FX�@:����M�����*X�8�A������YE�R\*�������M�N"�\�j����4q
�X�O,u/�N��м������'�{���v�Z���f8�Ԫʯj�d���(��A&�L�<�F����cE�_TQ0�7Z�����E�i�Ԏ�aTw�B=؟͋��8.���������VO�f��Z޸��ɜ�BV�G^xs��u�+�V�B�]iВ��.pN��!w�zѪ�{���N�u�j=��M(p;"��m�7V�и"��d��
�A3�V
'!��SNӭ�pگ��$�3�|�@�>%@̖���Os1;FT4pv���}�U��"P}�|��X�"ղ�[��P���£r{��/`vE�!�������Z��l|_�'�p��Z v���RQ޽bQ�CG�̙I�Lu1�x��Iڏ����q))���w��V�o�_��K6���@�����gØ�9j�i����%��C��N®�M�\�ͥI.]�t1���Y���}b���B��
&�?�5��,�WN�uoE���a�5CĴ�҈�E=���5��w��B>v�\��a"G�me�2_C�!�=���aI��PR�L���*������RO3����o1���:݌pT{��A��
Xj�]���.��1"A[�� }H�T���Z't��[X��Z��}��YL-����`��y0��p��F�te���(>��oZ�pX	�X�){�N�v�C�����#��)��f�=Y�3+�a����/P���d�uޚ
u@�tHB4Cb%(�}�V3B��Ѵ�h��� Vɂ|���^�j�n��Y3��6�ͽ˚ (bw�M����Jg"-`�ׯ�.��f'@!f���£�W'ogx�ZB_x��Z�r5|\r�{!|�zM��#P�����w�Ҏ	�n�pe�T":"*����9��3�>�Ì?��TAK���J�`�zz�
�!䕘B��b�7m�����p�X,#��L��d�5�="��˚��h��*�L{��PD��M�w�
�a��ȫ�\٣��uB���BZ�U��b��7	/����tKZ��eU.�a�Tg.��p�>8��h�3�0�Z"��-��V� ���1wU�+�-o�����뇦�,k'aHw�4a�a��sҌB'p��$�ʷ,���w�F�[�"�~m^"���>5V"��)�k��� ��ʼ��O���/�pD��;:��Va/zE�0_rKNu�%~)0�|�����]f#Z;!��i_^�oo�Abu�%�]�q��*��!);~[�J�Nk;c��"�a��Έ�f��5E��	˲%����I�lX��\ WS�g� %�C�B
*:�9�>���I�fx�iiQ���z�g.���%��[ÅC�'�
�¹^���d.���F}N�uH��ݬ	��?�aRn����J�5pW�fԡ��K$��ہ�:�Z��V�k��іH�c}��A���R�K(�l��&I�k�^8j�#x%\���7��	��C��m;�A[	��sĭ�)�5�����z9��i�Bo����v�+