XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����F��\���	CX5�ˁj�O��?R�3c�������� 
s��
žA�
h�LW���~O�&�=8%r�ޜ�k 0���vD�R�_���C2�eZ�N�\/�4n���&Jd��c�V��$����/M���qߠ�[fj���Q����PD�9g`=MqF��ͻ���0"Ӌ�Z�^tT4oj��7,��W�-[cE��sjNC-�ՙp�1�v1HT�&��U����U���6���F6��~�o	����uȏ�뚚>մWY�b�h�Ư����Z�*�|��'�4J��G�ϡ��m0
q�I����'U��Kb��Ăh;>�1p�5U�K~B��?G�mg�{n��\ܿ�>!^	]�#A���h����3��4�]�TR�p�:�'kY9�x!������A�_�3�$RE�� ��z�8�����W5��C+?%���Cm�Q�z���'ܤ�
.e(Ȅ��	�<��_E� ��$��躎�X��r���<��,�=��U؏� Z�r~)���Vn���O�k&�,^�g3�M�ȗ�/���F����7���wU�&v�Fj��NBP��T�����sXr.���M��Hl�;��+]<�1�e���/��:y߻�ΆdH�PYxS[���%� ������C3�JQV޶���RX����<×])��|
���T�A���풓3����T9Jd]_�&D���LX2SEd�U^�z�a�D\�BI��v�5/e���*�
`':˭��m���3�:/
n˅XlxVHYEB    fa00    26e0�Ja�;d�A]��qSscf��N��^�
E��A%���2{Z	�G'�2���a�M��s�j#,
)tj�"w�Ī?��]�U��e�I��
�ݻ���b Ծ�5��o�k�=!����������)��~��fj �C��2*�X�Oc�2���iCX懔��o+2ݙ5i*�9��i~���#�Y�X��}U���E�?_oE;�w ������.)�Y6	bK�K�{x� �|1V';Ap{p�2�������q��o��NO'u�:�o��I3{���K~�!������L=g+��/�槀�ޛ�֊ǆ��z~�Z�VF��
*����,���69�ohw��W���H2�/|�=nt��&J�3�ٙa���BX���]���9�?�zt�Vq����a'��=8�����4h�<��u�@��w�BY�$:�Z��-���0���Z�/�J\Ф���ԓu o��?R[r��oe4>kUR�wD��oxN���'JM������.�1�R�[�(��9"�z�T�p)B5�E(h }�~�@�l��G�J��eX ��MN f�xe7�l�͚�J�����u#�����$V�q隙�y�`�`�H�Cy��uR�R8��u���� 4 O	�11�Dƴ¡�H;����8n�k9�AF<U��`!"�N�`v�x@ ���0�;�C�>�]O���a͘�E�$�Wx�P���s��@��_��"�dp	 j�$���+�eb��2<v-�����}d�_�&ׇ�f>���ڇ.re�u	����ǄE�/�r.m�K,��Hp�K�pvWS�w���]?"oQ�&�ٛ�� h�`���mg>���IC&�ȓ\M��)hM T�>-���
�n䜸�W��	�N��	�gee�ʳ#�O�*�[��R�r�`�(��Ý0�7��W@��`J��e��?�fR��p�"  �=R����ѱ��LX�%��ٷ�F%�	A���y���q���]45�,�J�_p@�;	D�T�	k���y}�R孢Ξdޒht
lP��VW��u�{"l�!P�ޜ�vH�d�˦Q���ηd����!���4���2�v�QI���<ۛ�|���OOȗ�g2-l�J�Ɖ��X7���p�H���n��/���i�i^�%H�">X��*�X S�^��e
d��p�+S�,8>f���b-�-�@^���͜�b��+���^�),�B��#Nѹ�4�=��Ri����`�����35���O2ڸ����))�lƪr�t	w���5�Wm�L�X�!�?�����?�k�L��zE��l2�2�tm���˾�����Vԃ1V&����/ҥݨ,���ִ�E�V*�ʓc��S���j~էW�,�L��(w�T׷غ���������7��?,3�c�W}X�v�s�_.,��C�\�-���"	@�����!�k��>B�a�K��0;�d��ԏ`�K�5�;lYo���%ҙVۂ74�Fi�!��8�&��C|Ե��72Jkr�0
�i<duv�Qt������)���0�3����V,5?����� ��R�������o���I�9���w��Ia�uy��)l-2a���E%�$E�0�+�]4�����Vw�4��|!�b^�]i��_����`T����:KԶ��A����^m�]�'��̛�s����_������~��]�$������?�ia����T�	A�q�"8����lU̘'D�m�������&wO�GKPgQ׮�����M ¤G��rP'h� �(u���> g�]�
5m����x�΂�����R��S�]��\&�ڻ��,'����[C�m?��S���q$o�tx��{�o�X=Ԥ�oH�j�>�,.	��n"�uJd�3�&4��;q?��"6��S���{�5yFչ�8l�T�(d�)��J�t���W�5�޹�����)�Ǹ+ba��0Y�oCd�Z���O�������r0�{8�������ꥇ�Ӕ���f���5gV��X�
Y�2��S�m6����UQ�5[n~������3������D�=�#~�_r=��>-�-B�饴�����`��$�-�
�ǳ�/�Ԓ����Le#Z��-{����3�����ƅG�?����KUŞwS��� y�;v���=e%!o۪��9aͻ/�*P��2O�~�pC{�H�]۷u���,����U?�8dAn�Ȭ^�z�Q�0QG���y�^�z7A��JW!�����qV�M�[�'�X2���
�dI�����tO������:3�G��6;/K4�Ņh&5ę���L��!@�b�s�9�=��P(�,\y�T�Uۡ 6��]������I�Dl2��'�1̃TYur,fۘ���1�7J1ը��>W�����Y�93yQ��t..�T��6��ߓ孜A���Ѷ��0��|�Z���<�u��(�Iq"Φ���%V�T�ŌA��P1�''�{8F
J�SF
&;�w��8$�F��Vv�9a��.
�1T��!��9cr�S�#	����+IiNײb��PMR���NFܞu`�;	�b���c��i��Ǡ�������ޅ����o�?��W����3�Y�a���s���:ˏ�(��,/�Z�mԵ!]o��2mGa@C�3�4��$vn�0T���73p���(?�&]�����ST.�2'i\����Q/��h�h�H��G5��k�?�W��f�3k�lS�W&����3�,�����t�[�i��H���^��}��JRr��?<�]�q��W�6sޙ��O���~i�
uDD�zo��\����Y5kLo�� �+�vR�D�T� �''�a���^�}E�	Bĥ��`/M�����m�|���2�R�\Gyʨ!�.|r��]��j��zrp������A���-���KIl�*aW�zB1���W�y��W1?�]/L�+-������r��|�;���m��������BS��	�K�����q�Y�щSk^#�k�r1�o�Y�1�^�y x��x������Eeް�oCu��#/�"�]�-2s;^�Rx`<�V�o�,J$���̌<�d��.�ΐ�sC
cX�k�vkk�V��[�^�aթ��2�_^��.�#��O¿�h��1a�4�y�X�v[�LُY�d�V@ͣ�����:���~|�%���Г	�I5`b1+���=������D�1��'�ӧ��۽FH��c�ȩH�7���N��vU�(*
a	�_�?�;��8�3�6�$g��J4%�h���z��A��p��L�q7�&aY~˾�LZ~���*G�%�5R2�$KZ�hL��}H6_���MA4f�A �U9_�,4]��#�����0
�Q�!Y3�E޼zs6�H�.��!)���Zz�ɨe���P�
��#�Xy������,4����'��,�V6��Rc��Mfr���ݝ�{rT^�2�������<!�B5_xN~�9��4y	aD��͗G��ZP�3�hS��{_��!�
y��d�����L�uQژ�h%p}8!E�Y)�*�y�Og�^�$���8~O9C�	��;j)�ჽSl8�ܽm���W,{.�'zT��Ϡ���?��Xj����ڔI�Ros�������������Hn۪�H'E*�W
�G؁*�O�,a���8$��GH�v��.�BYM�G⡡��t�!Y0������X��>Sp	�^��ޢ^<����ǩ!6����J_|X]���?� vf$��5����U�K�C���1��#6�����ǚs�VaK�?�,��W�P�&,�;(�2�XI�gg�G6]������.y��O��ӿ8�UaHk��Dv5��@�mi�J������"n��#�J?��Y	e2ܹ����wG���:p,����ɧ-��"����O��#@���6��3��KH�!`[k��S��)/�g��nwsW LdL1�C<��?U��ʵ��+@&�+�A�+�^���D#��/���5�H�)5m��z�e����l�M�kノ�*D�E�!�'ꢬ#X~>$�}�!�7/]M=�h��g���w�+�����CD�|��`��-�h�*4O\���B[�ƨ����i���ˋ��������8V����h�jx��'5,3\��z:�Yy��^m� ��{F��*榃�JK��:#O#z�#�ʽR�/��p�v�/k�c �:6d�
�_����.�t�N���\z4P���c�Ws_�e��N���:���1����4���(X���ZtΦSz�fe��O���R��,�/J���p$5-��$U{`�ه �|��iڈ2�`/�#G�#�G���K9�w�z9�)4�?}Z�H�ݚm<������O�_y�F�},G�
�47�ȱÂy2���m����'�/��bP�|9��������p au�"�|�r���Ĵ�%m�`�;]�٦��͞�,Ӧ��Nv2s<��w[�+*�h ���5�2��)���p�x��D[��l�U�S/c.��~����'�@(�v�h���s�T�����JП�H�S_�s!z(�A��?N@�`d�r,U#��AYA����{�k2F<1�XLw/6��=�������Sߏ	�@Oi���OW�����Xc�pQi)l�C�I���ݟ˨��k��3 ����3mT�KG,_o��
)��zz��U��E�B��g2"�͆e��i߯��R��:y��}�̂�e,�{5"Ks00N��x����+�F�p��H�wJ)(���}Q~QkǓ��ub[�O^y�a:� ����ǟ+�]��k�C�Y- �f<� �����WjՑ��U|s�>��7�u�.j�\��Q���kx�Z�N��3lnd$CW'F�k���kH�*��VE�U-����M��:�rUe�d(�3���m,������j��ks���s�S��'D��5��)����M4�qUO�g��g��n��G���~��+���r+�w�ED{�۔����ܺ���� H]��Q8<�\K+?�Ր��M��s��j��0�1�Dc�O�P=�=9��jeU�-��JH���椐%�%�|Un����!��:8�>�~t��Ô0d_X�TB)�^�GLe1W����ɏ2�E��a��g�$��b_b��H����"l_IE�&&�φ+<�����o�,�g�v�x��[�)�q���v�<�����k}g�����?4���WT��+`:�P�G.ߍYDXܐ'6>�HrU�l�D���}2�k�<����<�3Ҵ�y��'e `��VT��<A��-�xz|o˂`��n�\u�#��,�����|૾]��Xp:5�]��f[�jxJxQ��y�%߫SI|�;5٫��d��B$��[�SsV��>�JQ��`� ��ђΔ�l\�&��g3�ܝ�����������A�ϰ� �;�E���o�HW����n�Dp�n�]�� 0K*.���c�X�%H�l7��$Oy׃�A���Ik~$�+r�Q$bi"� �r�Ss���Y��Bć9�֠x�\�;�~m����GC)xܡg+�3�L<�=�L�����!5?���~����qe�_�q���F�,料{�<�p��M�ꤡsA�Z c1o)Ŀ[�l�C	T�sz:�PZ_�B�@5��+��=�}n2�8;�1�Ǩ�qȼ|uB�@&Fm�����\��˱k,A��KP������!�ʜ�0��SDb����
�S�4�ƼW�k���,�;7�N�	Ti+�E��ĈTw"k�Z�1T�wмDD��<������I�w��[�p�َ�w���gh�ճ8D�:��l'R�ޑ��@.Q/:�qɶ/�iM�7̳/�:@��T)����J^:�7��#��umD�m]�2$��S�*(oa�p�Ѐ=��x]{�ʍ��am!����P>�m�I���Ki�vd@Ph,Z��p�DF�.�?�%$*��l*�:5��T�b��9{��%[�Z���K.�=L��(��U0�E��aO�|)B$�Y�!���F�����G��Й a��>"�w������k����Uj�]7`�Y����>^d�.Mh����ꠗd�%�[�c�0��^�a��.�-�%��J�E��B���@L�IO���6}T�xǼ>sPa�������Ȩ��qç<��S�)\tDj�Ղ��X9/���$M^]C?RO�UY��,!��E�*�,��@�%��Re6؝�D��V<
�j�@��Lu��F�l��!�t �B[����|z�����	�a�$�Q��Ď~�' L��o�ces���O��49̮����-�d��0����y���$˷�`�	�	�@� ��%��z�R	N�PDe�}4R���pD+)$�z�VxL��ڣx�10,�ŷ1��N@�D�Wۙ8j��KFe�i`�e.�~���	��q�jV�y�z���Q����eKa������i�����<���ל�O�d��L��V�:�-�� m~=��օ��B;^cS�,�u�)n���~��~����
���i�I�k��[��;�"`�ۜ�ZZ�U
��sL]5�Ғ��X��7����lo�m(u���|%���1�IM�@b��w�	��ObU-
�v����T�f[9>����u��ʵT�:���v2�E8�-��Rhl�ڈ� ���q !P(qM��`7��:S���1Ρ�J���1zli����"N��JB�}^d������Q��L�$��c$H|�Foב���m���k�*�
}<�|}�W-ߊ)�������RRS�m�p��#%����ɵ����WƜ�X�;�6c�/�ֿ�\�'�/� ��)������]�I�9�Zk�6�K�r���Ѐ�:;k�ْP�0X$����<g��n���2!��fP�'Ɍ��b�0_954��?��"&r�3����T�4s��g�@L�Qk�jK6�
�]G��/I|��nѫf"�P���"ؑ������)"9��v��Iw:�Sa�P��A9�eܺ����?/y��ډaD4 ^-O���UC��|U��Y��h�c/0P��F���lЏ�p�O�ѵ�l��
wp,gÅ��E�qhPN�U���͛��5��3w�k����;Y�|e:�̰]`㿟>}Z�5E�Ou�5����q��iWǃw���J�-�E
�+�+9$���F�#-�Ƈ@>���*y[W��6�d���4 ��(�2�2��Q?�2��u,r![��P�����A)
�f�s���(V��A�Dk1hk�l�&6zSe��9������%覔��?lh�:�����)�g���x����$4�[[�t�|	��W��U���K���[�r��qW2�:����w��z1%<U�JOt��tH%��[,�a����:	�X���a�֯����n��]�C�?��"��Rx+hZ.�R�r���~�W��� �;I��������"cr����cmM���⠕Ƚ!�"*�|�v���V�'9��F�P<S�]z����|�R�`Y�";�fU���r0Е j��&javq,����\&bo�y��6��db����%���MR���ܕ^�%�Lev%ex_� xx��>���i�x �m��9�\Yt�OdF:�aH���!���Ǹ�RI��U���7ᘴ7	vU������|X��""*�_y�tډ��^#QJ|����Fi�쥒�3�"E�ù7��0Ǣ.3��Uf@��@�*KL�$���[�ė�AG��Z*��L��c7�#=F�J�U���Q��Z1Z���Pw�"p���t�{R
�R=���T�vZ��׏m(:4U��}�R��N__�Ц<�r� B�E�z�¸�m�����|':�����.Z�Z(طj@�B�����Q�r�3>|��m�5L��$B���G�C��T�:?�!IJ�)� �-��9ֵ��۶ qBB��w͇{���خ~��9���IP���DXa��r��s�(�A��o7���=P_��+>ô�����%V1�UL�k�?_
-g�Z���l��ی*i%|���fn ��;�?��C�w���,�B������T��T%h�O���Ɂ!�����&�F�����?��a�WN�t�����0�ʨu�����5eR�]ܸ��04}k�G`W)P�\o��f�)��C��2h���R�a���!�Q���i���ڦQ� �R���*���e��y;�OQb�5�1T����ZLك7՘���O͢s<��w�,��-6A�Ԡa����� }���Fi���ŞS���û�����P��B_	ng|*���M�l6�$0�}K!(Zo�����g	�LɃ$��X��;4�[%Z
S�"��Rd��^����>)gL�9%"���C]���W�?�r�\o�&^,H;m��Me�m�g-t^�&�IA���O��4��z=�3)m��AY�}(�4|Z�ׂ�Lr�Aq<M)��7�5�S5'�	m��9�g�WWI�/k�E|Z@G��)�9LDc��䓵��;��}q�"
�1��?�#颁�,��O���E"�?^�4�՗<��na[B���ܟ�C�.8k�Vgr6�� �=,$G��dd��?u�I�U4/U�+���r~.�$;�t.��`�l0���`u���Y�����+����da�2YR�c��2D�	G��Y�Z-޿ɾ����{8��[5�w�3���������1{=d-�'jl��?�J�8����9:7�Y9������U�� �9J�g4toK 4��|�.US8�m8]� ���9]�E����(��&�li���!U>/z�9+�3`�#{�z.�eDܽ��:hᓹ�c}wԠE�f_='���f5u�5��gcJ�6��� L��|5Ca�[K���~���'~�v>`�7�<?��5�ɗf�Ʌ�\时���:+wA�� ��C��Ɣ�w���v��b�@bs�KC���+�,��$��kq��P�oo��$�nQ}���U�8�h�j��x�&���&g`&��xj �ߘk�#�5��Kyz��s#��(�����i���M�
34�� �k~��+bd��\��S(����Z�l�c}�[��yu�}U��y���x�4�@/�\x�}Ђ�^R�!w�f���M�^���	ZԨxA�q�Ի#ph��/�0]�X�!����z��z,���|#_Q�I���u��0��H���{�v�i?���vI�� Zx�1n�s7�a��BXׯ���TkT�@+J_� W,vo�k�����yN�=_��?Zm'��FSX@:���k!��s���&6g��. ��Y�
���[3��5筺c�>�;49���%$^��!u7��_�2�6��;:�6����6���H���/y�X9)�)_��#"U��$�����a!�b?r3m��g��Ίկ����O��9�Q�;>=Uk��҆CaK� �����g73��E�.�F63�U�z�Ț!g�V}ɔ�"�$��7Nga =l�b�yQBdX/���|9��Kح�vkt���������d�[!oA�e�Hv�~/��4�b�����_�m�NG8��z$N��/���p	�t�
�34m����&�@�#,{C��_�<�ٟV�An�	0�<���D�mRik!�����#�֨GZWM_��]Ð�����R**������>�$�Zd�r����H���G���T��a�{�����(�xA���r2o0
�L�g��"��8�b7�߃����C7�)Z�Ɏ)x��̩4r�9�6Z��Õ>0'9+�f�p������m��"��"�:^��3��C�`I��!���XlxVHYEB    7d55    1450�^ @Bؔ�Y����L���P���{��N�+?�Ae�21e|��
RQL�`54ݬ��J$�=�4���#Ǐ p�BZJ��^�v�	�􉎄�^�e�A�9 S��]��42C��K�@b� S�z����� o�!�;o���Z?��7�K�H����U��u%�� -L�䍓����v��t���k�� �|����G=�:te�q7�w�Qy�ֿ#Q��Oڍ����z��m��k(��S?������k{N�����A\T�+.BZ*i��~W�HM��i��B֔fdC~�6^�)����=K�06����}��@+fc�c�C3�� y����Qa'���z��2��u��I3,`<b�1���)�&��<X����ȉp�����R�*Ԧ�D^��z���*|��1��,D�.�D ��u��Z"�"�����Cg�0{ؼ�`���� �WxTb=02��G;V)+}�TZ�Ns�r�EK�*�!z���6��7���' L��#�^f��p(4 ѻp6,�~W�y�c��xW�SJ��t��HH�J��W�*v���d*\K��Y˙�	%�Ϗ�+Y���8�;�P������4�ܻP���o���E_�]�5ƥ~K����ھ�rV��m8���������W'�O]��0Ɔ�4+�-Y��+	Q�2�t�i�͉�ǹ��uN�oɲ�ԯzM�9���ld��X���桦q���|gE����=.�V��ρJ�Fy�*O"V@��F��G/�;�m���K�"X^�e�����m�C���񆔦���骩�*j{Nu��̀�+��&/1%i`O=��J�x�!�R�ԕh4UH��|d�bh�?z���[�$�����
E�n��"A�}�Ӱ*��:�T��h���(/4/��E�1ے�*�6H$Rg�g^�C]{^n!S<kO��
8�bD�"96�j;[I�m�@?��+}Uh�,;���MK$����c�פ>����(�Wl�h
��d�$E�.p��� gw�W����ub�E��J<)ty�>F��1:XR��aF��Pr���/�Y�]�Up��j<�s��3?[����Z��m��9xH)�&d���-��^�z���+�f\��I3Pq�pT�CS/�,!�\�-h��43uK;N��\�7I����q{�v0%��s�B$�O-����k�m����l8Υ���r�k}������Ӳ-��gh%����:�X$,��a�kՅs�yxWC�!�%�gk�.y��;jd^��f�,��g���X���
C�w��$m��x���?��lre4��4tP�`��T�I�-�WUS�g=�`��H�ސ�c>P����ӏ���t.��[�<�㲀��$-�>q���k�Y,nx�D7���[D�ew�s�j¼�
5c�x�����^���3L���p"�����K�����c2�?o��v�p���ƙ=�)�K`��̔Sc����5����]^��x��`S��Z�$M��Ƞ��G��m�{"�L5~ar�W^��W[��,%i\�)�q�������#��
�p0��3J��t��x�i�3�q��/:n��w���^�j��;����O ��2�b�� ��Ξ��>̂��{n��H���6���ż33OTQ�0�c���+>k��p�j�{-$��7�Lt[ۖ�%�"����bm��:*w����.������c~z���^�|�ʄ�q�mٽ�K{��`l����rm��L��\���7�2,��3��w0�&�J�_R�MSJ���䐩E��<�M���Ի+(�Y�`��9�R�6�+ S�ꦠ*���{a�Z���)�j�U4Q9��F ���]q)�e5i�TvF�Sb$)@���7�<�(_y��u���_������Jo@}�Gˌ��1�l&�Yσ��K䧝���1l�_t��(�E���$��U-�hX&�OX�w���9Ӗ�|{�W�
�"�� b����Lŋ�A��)j�����ht	0e��詨Ø�����֪�qp"��
�[_�����6�/�W����x��^Ej{4Ԫ.�E�q� �KE��WT��,�BZw�-ɦZ�J��UT��U�<�o�x�	����v��Ă!�օ��J���.����"SnIBqC�#�����:�mtj�J���e��A1�Mc�*�RA�˽9���co��a0�ľ�֚Z�L�G�T���O>$�(����+]�l|3��p�;7Qj�J�B�f��sK�gp�����3Ʉoh�Ft��I�To�zT�d�m�*-gg�#��%����m�U�ϥ#(�KS����?;�B�#ް(��D%4>r?�A�a+�-�D��.!zSK��⒂X�g��B	� �jC�W�p}�U��;z5|���4,�WM;
��N��M�Vv( �o�(����8����2����q���`G����B5Hh>M���9�c}�:Ŝ��,?=liz ��Λ�M�I|�郪���lP�����F�%�0~C�/7Y�iצ�e&�_j^�lJ�]!,��bwg�t��h���NlZ�R!w�#FU+�$N����%{�x����fÁ�n)���Ҥl$�h;:!�[+7����X����!ֽ�T��Rt �{
��E�O�� ��ϱ�<B�-£� +��<
�TƔ]�R�o�h��jL �Ob���N��2η%P*�ۨ���d�ߥD�;h�z��-+�2&�Q[�v�����Xq�������>-('�/@'��W����Ft�0W��
����ò�T$�Tu$k2�x���P��F�8����V�M�^w-��|LN�lts�ß�h���j��N_w�I�{T>�Q6�j��X]����
f�!�p��=���x��r�ݥQG�+Ń`�B��5	.�?���DS�L������!b2F]��6
���4<evэs�:v�Z�$iB���k��!�j��]ӥ����[I�b���D��Jp�Rg��j6FI&]�z�mGy�I�cr�|{N}E~9Q*p�F�n<7w�*A�9���>�����ݫe��T>����8��ب}aV��b%fkK	����=�L��3!�X�M�rÂf�d0]��nj 	�2i_Ѿ�x��7�k�I	��{5L|W�?�h�c�pL�ڗO3�J���Qt�%��+�}�oǻQ�o�Eh׳%�<w�}_�����@��ʦw�w.����7#%�T�G�L�s�M�������?�=RB>{�u1�_'�8��FE�prpnQ��-@ ����)hdVk��}�n��R5�$ihlj��J�������
z��
l��4䷃bA�M�J�S�� ��ӨXT�P,�
���_t]�m��|�K3|*�yE��:�,ĒgN�C##z�^]D�v�bW�T1�1�I���ל���=_6T���?99,
�َ�<T������X|r�=5_F.�$`�N�?���a ���00���0&���)�i��HeT*���hɅ}�Q�q�Qb��wp���ts�6���K��8�f��˹���u�Q�I�ˬ=P�Z�Ҽ�T��ed��O;�.�|�	��&E^Z�RY��M�˲���]���e�VU|�T�u㪛�p2�r)���$81VF��~���$���?��FK<Ld �;�l'��<g�Ȝ[���9.�U�J$�o�� �V��p:�u�6��Gf	3�OU�X��\2�����T�/?x�]o�q�=%v� 3����͸h��%�pV�c�,��$d!Dn>��=���/�Si�1��jl���#�Qfq�Q��h"��h�jĉ��v��^*��l�a�� �~.�]r)���5��ʚ�i����`��s�5Y�j�(rX��δ�n`N(,Ҙ�����G�����:ލ�cߎ�r�"�l����5���]��{�mW��~G�3��Dy�e۠Nn8�
��fr�BxA}�4�-�H�pz	�#��ac�����߉�E�s�LM
�<� L�)�~��!X�R�����*�2��.vA^��=F��sU����,X�(�O���x��킁��
)Y��Û��%/DH,(j�CLW��ᩚo%���(����ЅȰX�Bd�[�Ȅ�R��:�BΡ�sO�
��׷%�PiM���9�w�����M��X�e	5�KF����_>gc�?�"vb�A���Sw	����&,�#�?�(Ƶ�g17�G��e!��n�G[,�W_G�K݌Id�C��$rU���%�y��-Ā�i�S?�7.�D�Ik���c�9��69��³3�}7����n[-T�#q�b�v�q�3�Å$uξ�>����l������E=�Px����>]X��������l�U4��K�����@�8�̾�bS0�J�*���8�%L�A�V��ښGh�Zzs^��C[��XG1�c�F1�O�1z5t2��U������,�q"Y��I�AL�{G����p�Rۙ*��0�x6�Z��ޅ��_ "ZH������0�iGGr�����.*�fT�K5ׇ��8n�f�n����E���Y�}���3�?ɟź�P�<(5"C� � =��
1ؠ
��Eq��H�����J!S���n_V5���3n�~�y�Y������#V7��t{�r���P8w�r��6]�t7�Q����G�z�b-A\��%ԳL�3G<�Ѵ����_p����Mɤ�N�W�j�j���}?	,Q���+2R�ځ6����,,X��l�4LC�����88]�W���f9��f}+�ǝ�|�����o���*%�z(�:�j�����37!g�*`����n^q��Q��+�Õ$�IUcL�u*S#�@�A8��U�Y�8��`��0N�9�b��)�	�<Z3��1A��Q�Fk`{6�kYc ����v�:<x(0G�O<���¸�X���'XPXh	�������b�$�I0�rZ ��w� ��;W[�I#�d7]����8ܢ�9��l��?�K}@�l$f[bYyDK#�������|H��P�t;U>)�?���ȏp:I�%M��0;q��Z5i��]k$� �$��('M��cGܣ�(��o�)����(i�S�����5��zYf�O�N�'-�Ѣ�*�#��L"u������|���?�X�_�C�݉��C}��P��
M�Z�K��#��4�XV��