XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���hXX���[��b�څ5��ڞ/�L���J�{x�t�h�C���4�:��أl�'��`���'w�9��./d�6�lT�?>���=���%Ai��}#:���@�#K"K���!d�9�b�vwJUu�\y��
�U�����9x�h���7dR0��L<1�|�?�M�c|�=|��W1�GAD��X��ɰR5I��Qq�jFU���^�覧2-�[S��F���3T/QT�����[Gy4Q'����V{�fn	���+�pfZ�`1�+�ږ	��O{��s��w��َ�����J�(�'MxP�*�>��>����p�� P�gQ����)X��7n�n��W۞����S��[�����̋�^�Os5Rhw�~9b�vG��<(\���.���칱Fc-5 YC�0mە��C���F��G/�ϊ��8�r*ĥ%s��m�t���X�gn'*y�n^I���T�;_6��y�dp�&T���Z���|���5�l}�/�{7:�h<n��;,g�4p�DH���j4�x�7)�3��~Az���)��ݱ:��s-�~ε��/����]�������[���w�ԧ�;���yn�2�D�P)���:j��a��$��X=��sY��v{+J"��W�7�7:��,�]s���g{w_�`J��#����c��wмjnh�K�N�������?1����Ztg�>xUl�c�jْ-��!q�Be�L90�"F��wA�V�� 
v���
}u��_PM-\�*���n�O
�u�XlxVHYEB    b087    2540��,zs��~�u�S噌2�����a:�pmv�[	�Dq~o�T�4�%}����(�T�����}R�~a�-���3B��׹< ������U�S�\B��<��s�}Q�c �m\�F�~N���Q,Hw&U"M��g���昅�D�8R^u�M2l�Gw�)�	���`C���6�7���	<|�%��5RB��-��Ԇ�+FB�jc$?�@��h1��3����zU��h��'!� �n\)�\,e�HUO)Xe2�LܸSL�ۀ������U�q����] a�-S�.W"�Z�G�=r�� ԭ�te)�$��zihW�TB_����3>�D��{P2�D��f��5�~>CU	zL�
��~x��[����v��i~;����)qF�'\{���b �7��Kt:ki��&���A?��EOj#Ġ(��BĂ�(@'Upc����LХ:�C�ג	?�g���I5�:YY��8S�n�ci�_���<������c���9�=m��oS4��H�M��0��m���}�Q_�'�\V���X�Ș��VǼ����N�#(;��@g$RQ�1֤��=�O�Fo�M�k�"`8�ԑp`�F�h��d��j��$mr'B}��\�ܒ���$�{�?���u�[�Ά�,�xn7p��I��2i.�ʝh�ۨ<,���	��E���]t�*�PPS|���ќx],}�#ځ�T��M����A�)܋�`�UTŖ7H;DV1#;�/����'�Hd�ğ\7�LR��[�q����e���R�~�)Dpp�t�JO�h��d��1*�c@���퍋ͦ���Jd�Y���K����GM%��]}hө��*5�Mb���u��m�_Kt~��I�v������AO2�jM�o�%��(�	�^&����#��)�j�,E��ˠ��8k��)J��n��[����=�x�-'<�ڛ5�x�̾��Xf�cU�~p$R[�J�p�<��D���w(��;�G�f�������ǌG�L�n^���_L�*=n&G�3��_:�-�qhZ���{���z���)��~
K��#�-��;�f,M�a��ڨ--�W�
�|�+�i���9�b}�&e(��k�1^�c[]A�T^�$c��t��h���v(" ���&,�d���`H��~�K��	�4^/�g��H�b>V�B~��=�����%��5t��TXJ���#����:V�NT��M��`�e�哵�G��G��f.�^H�QN�z��6�".:]M�E��~?>͜X�KQ��*��Q=R�8O�Te$ ���^�+2i�����YǪ]>7B$��s�bDB�����W'�z'ػ���l�E���}t<����T�N�*�j}(��'P 0���z@�N�XflԂ)��BU�\ݰ����Zn�|!�����N������h.P��#ִƳ>θH��C����m�fh=ʞ�#���I;Ӹ�}��Lc�,�[�F�Ǒf�,�_T&X��5�7��bq�Q@�U�sE�B�~�ѭ'ݤm�ʤ0�x��1����|B@d��J���B7Q��yH� �ۂ�b�{]�Y9	�!Ή�_�f~:v�am՟�(��غM�Rǋ��B�`�Gv�ڹ�uzy���0Zc�x��M-���0��K%�W9��l��\Y��S�/<��S��dOc��j)(�5M�r[/���5��/^NJ_����uC�!d"��庱��7�n��$k�-��U��P�&NUB��и-���پL=�ړ��Q{P��4���21��Fb+盅K�6�ٳ��>�XW�mo��l񣑎`�U�-� H�=S1�A��:�1�KU��pY0���%�w���"܈���VP�z;v�rn�Z5��o��e��X�`ʘ~���2�oAU���LS���l�j'<-ᨽ<��xfN���6�fl|�Q=�hۺZ\4�G������	՜f�����ް��sGP�2��RFq����f{I�V����l�	���L�J(;�c�s'�0��p-��On�q��5��J���X"m�\c�i&5�&2=�H��[w�L����R�c�vsE�F��{2�,ka�rm|4XX�m�% ���#�Ҳ�M,�FưP��Ɯ�y,��zw��<�έ�.W�u�z�>U��Nε�S<�z`}�����73��A1�<�W�=����C��h����y�w�����Z�K��eD6O3GS�
�3wG�Ω#z�x���n�TW+��ȏH�[��_9w˹`4^��Cd�C���؀}�k�k3��%��Y�r�'V�W���E{k&Wo`�zRtK����3Ҡwz��FM���x��]�q����֟E��y޽s�p�����#H�V���NnE�ʚȜ�������Tw7gn���{T����Rw�2���E*Aqv��ߵf�h�i�b(ĩ	��Vr�+j�;S���eWC���=s&�::�#��V�P%&v�'(�&�w;�$�X�7D��F�j�sCW�JV5�%�ӚO� ��x��C��7�� e'yV��ת&D���0)8j�K�A{�:5�2+͸�Ѱ3�ם����+�Z�c:g�	�tΉ�� 􁮿� �0� �����QG@��68N�K��n�υq��`�"1��?�9ot��./�-��Vt�g��L8�DFsؙs�LϜ�1��J��p����6�>�N���i[�5!�B����M�O��2}��TMV��1ydQ*:)�ۆ+߾��mUGA,I����"����k�/D����4s_�;	'W��*qDᮥɊlr[`􄤔�*�����8�ٍ��eN�+�ו�	�P��*!��PH-u�b���&�E;�y�!+�Q�\l\vK1�o�t����َ��\�� �5<�|��>�vh6���o8�B3�	ᾄL;�a	W�x����Ll�#����tX5��Wӝ t��2\@�<���c<5��&��BN��\f5o2;�C>g m��)fPyq���1'+#p��J�s���*ޓ�_��~�����)�:�dIv(N��������C��ō	���n�궫0E)]zC1�������q%s��E�?�Q�{>&��ݵI��G�B�ّ���J#�@���!\S��:<jGl��L��<y*~�_M0�,ЖT	��<���.;������q�����R�+���-���[1{�{Fz�N��`��q�t����MĹVkβ�jgQ���R��I�Br�pm�(�Оp���+@Uoܽӝ��?c-�V�r��ּ���3��W͆���#^_�@��OM�~�<K#M��gq]>aE׿-x���(�p��z��x���(�hGo���;�=e���ID�̯��= ���I�B̬^�  
�`�;B���8P��ƙbd�5�"����d���R9�ń �mZ(rT�:���xl;ׯ����YO��ǆ�Cc�� =ܜ6(#_~q
�Hg1SN����>:1���<nK�^�(d�4��Ô�+LK�-|^	Qȫ(�I�\��]�w���\@~��+�@	2ڊ,Ͼ���ٗ�6���ڐX���p�	)#��V>)3�+�:E���(���B���Q���s��+"8���,�G��ޘ��擟@�i9�A�՞r�Bڄ���M�#Qe{���hmH�"�6��UC#c���~$'�ֲX�a]��Fd,������#%tw�>Y��OF�H��^���X@t��.{]#�|�F��@P�����GXj��0�D�x ���c�`+�7��#DcObw�(&S�z���؞T� ,��b. 	I���v)ˁ��/vk��'�����CJ=r�u�=�i�� KC,ZP��{'�1�3��
�ס`��Wj���=��KZ.�w�D��l{��JzUϢ�;�c[�^2g'��QYC�U��)�92�(!�A�� ��xS�&{�Q�����Qm�װ7�.�߾WH��s���eꗅ"40O��2�ZA�a����s��a��uD�F�%�d�4�x�Y?���w��+R�ب��NQO*��	��K�F��No<�����O�sy�-(U�C�j	w��(�V훕[ov ,�������|����m���(��^h�H���>����@͡�]��Sa+8gAK�q�Iy98ah
|V�&�vؓ=ohW��������4y��v`��c񋾄SwtX�Ȟq���{0����H�΅0�0��oP¨hN˻Z�hQS���<�Ԓ[�&H�I�L�?��j���y�$��<��}�*�����*k��'IDTpf���V����,Jb�������҃��ÇB7U�~�������Qd�}Gu��bZ��
�дJ���K�j��ɛ��<�ˮ��?m��,ІQ&���Xe���D�s��<��u�x�G.AD�!�h.�
��͕b��cc�>�@l]lh�:v�6��~��x�>���n�D�d�X����t`�>�Ȏ�.uTGD)�}u(��ȶ=�����Z5�|�,��b
Q�p�3'X��o5>���q�{!�\Zu��{N���5���S��-���� �((��a�Mã�Ǧ���7���<:�F� ��Њ\��'s�a��l�-3>"3�Y���vl�7H_>Uq`������'��d٦�c�%O7Ƒ��:'��8j��:�������%`�.o��EZF
{-۴J	�����E�y�,I�v�
#�M��<��\<�<�"�k�wrN_�2�oY,D�i�o2�TZB|Sif��)\�ifN�YPwJ'�R�Q�Wkw�lR�.�`�/�m(y�W14z���O]�*�I/�����"RZ�}t�T�k '�P��a������A��
 kBf��_�{)�����O���# ���li�E�c�z��ky2�kzص���jEd8�j��|q�-j+�ڻ�R�F���<QǸ 6qW�w3��7b��P���"~�}��2����xf�Msw��2\{N��S5�KC�fB!g�0IQ6�C�����M�� �WB˳�l���"�g�a�`����A@k3$����Dz8���ų�t8�(ue��%0���;�0�z��l��&�HV���`oO��rt�H��d�>IO��j�Ud�F)�8�:����fY�8��l��UkF"�d����z��&�uX�j���Z,��$_���R�F�ڽ� c���J�ڴ(B���~J�B�H��@ɴ�d��,S��P#�5(R����/`��������s�����E#��'���~�{�����X��xk{w6w�lM�-@Ѿ���s�fN�s��M�n��s���p�ø���@̖�X���G����~o^x�
�&d��a�n�h��� A���R<�X�XW�Dtw0Fj3��`;Gf�	����z��	����,*�۟k�G	�̼%���i��/�π� I����P"���W-���e8!$��k8uÖLH��p�+�).=��}��N��H¤���N@�f�=TTs���h����̸�1K��QN,h�s�<�(h���.'?=|��Y$�q<~yX�������v��K�[G�UP;���4+[3S�{#�rQ�*���:M�Z�,��Ȋ/�'>9���U �Bf��O��s���ݻß^���d�O��-bfx|㭸�u��:d応lΩ���+�<�e�q��T��qx�����-f2s��?f��To�F�\���୺8�Z������:k��SF�#��;�� �6t΢��1��.��] ��h�y���n~��O�e?��k�y�*)rK��~�sV7���f�$ď!`�Ue�!Y�w��J9��	�@]AE��� ��]h��3Zm��}D��G.���A�_�W֗xUYz˹ +b�	�ò���ߦΕ� �D��
}֯	H0���ϜD�ʥa|����KsLC���(��F�Jɬ�xo��u��Ȑ��y�F�����U�VO�X��&_cԄu�fY���T�U=��ʘL��x� n���o�{�#�zx*O{��t8�����Yz>c��E�d�x =P�$(�z�����w_���װW`&�K|�˿v�Œ��w,T�u>|R.�cJ���ԇ��R�U��i�d���/���z+|(	����`8�!Ƕ�o�����_��K'�����HK�F��=2���qcg�LƞZq��ם�J�<��[��xU(N�n��I;�A9U��(ʨ(&��Չ�l�Sn(VuV��~=�	�7'������?���?ҀYZCh3��y#���O��<.�y}m\�H�"ؕ�f��G�;��D��{�>�U��9%�Ǡ���Bl�Y�r�6
�9��c�.55Cl�|H�����D�T��E�2��ƞĵ��G��H�5Q/}?��W�k�n�R㛐l%�cw��K#��Su���i�E6Ȭt�[!��>��1�H�t����+��p_N�Y����I��6��X�
�D�ө^�f�|���]�ĘP�V3М� �=9��&YL�"�skM܍���}%�`��Az��O��YC��߾%m�f"�ӟ��G�L�Ӆ�z�����@V.@��/����_��V{��qz*�Q�cn�%���hTtMk�lP��B$@�/csiNK]��s"��GQ������u�:>ux�G�As�'
�l8���ǭD$���o�:w+�zH��ȕI�n) l~����e8y`��m+�Xg�&F��;Ї��n����6qm��̄��X؇aqS��&Ƣ�_vO�1��N1�T�mp�!��ѿ��q}��so.~OE�QT.[��H��g�j��<�E�|��������P��4]m�(	�#
������9n���,�;�&�#�!|Ķ�\5jͷ�,s��vG���FeEkC�ȱ��ma[��d�Svh���_�l!��G�U��Ƥ��U$�Յ�g�D�n�J�!l_I
H�9�I7�:�2H�|��c�؞���HC�����a�n����쐭�w�c��
��U�/0����A����M����O5
��bk����?�>�!ojn�>��D�.�bu5g�Ӆ}Ka�^�M���'*�2�2H(�!:x��`�`��\����4�I���]s\�&W���No�)��IX�7!�l��`�����R�����W��v�S�,e��	�is�r�b�����Ml����.� ��� �$���+���V��[+��g?	!dg�~2�� ��x"�چJ����۲m��x�4�)�8<����'/�����*�߫�g�\	��}y���R�a�*N��x���@m�H�G،�IPe�%g��|�2�~C�1���V��v����[	������%D��C �;�0�����ZG�@�Y�k(�#���U�,*G�ݻlr%��n���=���F����U`h�~>����yI.����;�b���7��,-�V^��9�	�9���3�۶���hxr�(���*�m�^&O�!�8�8
M�T��b���9������a� �����乌�,4#�ן��_Q�b�����3-�؂P�5RU��qM�^��a|�>�^3*�����u��M�)gw�`(A;?ǳ�]������W1�R!T/����ñ#����7{�o1�Q�NgG�8!�;Ō�:�?��ՈE��+�#S����8���ѿ�lӡ"�^o���w7�,`������M�A�6�����[�����d����&�k���d����ZO���O�-�;o[��yqv0�#�d�GC�ۑ�\6/\,E�P��u:�L&C�EO�I��NU���#` �Ϲ9J��XOE�����8$
X��y��V;KCr�))��T�G$i����E��8y]T��̃�d��0��V���u�b�=cY��$_�8��1hΕK��+- �du���qn`���WF[�s!���M�}��_h�x�+��O��h�N��E�Q��t�-3��%W�㶤�w;�v�/3-�a|� �A��[v���dVի�!:�)�\V�KP������Q/���Կڨx��X�8k9)�[nsJE]7�!t��W�(O)���G;��u�s1/��&	��PG�ے�� �R������"O�Al
�&�JZiF�]xI�_|���~د*�'�Ӂhu��I�I�0W��'��U����;K��(�n9�7?^-��Kߕ��ʈ��bKf�Z	1_JzZeO�b)��_~f��R����%}����lh��x�Y�`�6�,���������bӾ�rbq��'�%���(~�]��5���&����%~�];l�����"F���Q��(ݤ�qx"��:M����������Ę��YkWMl�z5����>l�Y!�3���[�S���3�E�h5z�>e��i~=q���Ӡsr�1�V���R�摓"5�3���h��;��|�35�ty��B�J�O�E�yFH�@R��?�rb��
N־�v�R���='��A�P5�9�a!sяK���$�
�0ق�,�����2��dIR�zV���|P�mḏ<��֭�C���:Y
J� ����&��]X��pxj��/��|�&�t�;��o�b�C�n�v�T`�JT�]lB4;�?��%=�ݭғ��{���¬����6��,�7N�5�JW�AK��d�o"��g۴]1��'a���&���	��߃銪j6��X�?0L�����%��#z��fU�٥�����g���gI��Ch�Y��6�.�[CU���T�9"PFh��'�Ue��ۀ��?���K)�x�����o�/Ea~���Y٭��q��R�M�`_:
'�r��d�Pg���e�0f�^e�����-�P�Bĺ���}��)�cG,
Snِ����r9�s!.3�r����#�sw��!�}΅}j���o��6�w:�g��H��''�ne��3>�8���aG�w������Ջ�@A���$/R#�'�/�S gc��>=ZQr��H��*.�����gB�U�����ܢ��B.�@��\�0��
T;E��/���')�4�n�g��>c�Nݥ7��^*�+�	�v�<��w-w��7?�����(}�R�a�Ə"��
��=�jĔ��愾�v#L`�\�f�l��+"��j����Կ�~�4����je����=��9H�,T��r��zI��0����Ӥ,ȭ����۵�5=��x@l��ǹS�l�} �u^҉M�K!�����]�WR�a�H(Z��Q�Z���waF�<E]�u��9�dbF�M5�B�PS,$��e7	��>k�p%���+��R��On% ;�d#�а�l0w�,���6%���}�
�`b��o��7�}�J�6�L�Q���0��/��.��$�F�B���Y�s�zf�h�����^��4��HV�0��'T�ܐ�|B�ȅRHE��PZ+�Gzԝp���8�T$����%r1s�q��aI_�?u�sZ5