XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���q�Sb����נ\�\~$:M�I�&JK߱&��k�� �8�3+�Ǳ�F�a�p"{�K�y�Yl�L/_o�x��h��I�R権�nOq0n���X�X]�����*Iڻ�;!�c�%YQ6g�(�a%nf�0�f���}\a�zR%�G��/f���5�W2�0������ �K�!+F���X��=���#����P��M��Ţp~d�X�v��@Uw�����ٙ��y�H�`�{(�U3K���e.q�%��d���Ei+�Ն'm~����ˉ�.�Q��FI�n
�b>�9�F�J�<���j� ���~=L?�����-�=��UV��o���W���j��pv�YX��A�6<NZsְ��y��J��ʔy��2���0�l��a;�by$���=9D7�T�&�
�޶}U��ٝq��0PU�2ɶ�;S3�J<j���d����=�֊b1�P�����Y-|��}�~�6���#P߻D'�}�*5��a�z�3�G��������<k)1�8�� �X`4x�8��t���q��NB���F���-��aAGYXGS�nR���p��aYm�Ӟ�wB��.Ӻ8��Q�� -���&߾��	!b�!۔�3��fG�C�)ݑN�S���9�t�-��K*T��e�k��ٹy��ĸi�� W��2��E�[�Y�d���d�SGm�X7�)(䶥�e��20���@obvB���I#�����'�Ɠ���5���2��{{G5�l<WfS�@�1XlxVHYEB    6315    1790�� ���cs{�!�ҋ�J|F��a#��|��t���9�Ati�;�P�Ng�	�K�)tY"5��˓D�r����uQ]��o���OYL��mx3����3@��D�9����;��"�.N����D�|�,\� �?A��|R������ɐ�ͮD�dĹ;|�cݘ�.���A^���
!���[<ʟƚ�_+��°�@$[�l�h�h̭͢g��l�ޡi���8qt|�D���;XݑN'�]ɞ�k�D�
��'~��;�*��Y������@.�&:��l�)�Q��g�a���a%���a�Ե��4BX� ��$G1������;�Rt.g����(��9ۻ��Ĥ�1�Y��(��>u?t��۵|&yk����㠡�D0R��\��:Ѯ��-�j��f����>�։���
' D�ȫ�E����=0������R�REah�P�I�`�拭�*�h:b��Mo�a�=��?�P�����;��^+
�7� ���!m�W'iZy�<Y�G��a��!�aA��v���� �����sAa�s���w|ҽ��݉[Q�e4���P��Z�=ɫ�m�mV�*8��%��|Ҁ?of$�k�4�";�/���>�I���](�K(D­�KϔQ�ꚬ��|��E\�:=;�?�^xB�>�y1-S����VDE������xʭ��5�G0q�Plf,�2YM
���b�V��8�J�%'ϓq:����%K����O�`��n	s{V�Q�I�iA��I�����b�S� S��sS�Ɵ����"��f��ի�7���ۂqq����O$U��}{�S<=~��O��\_�*e\UͻG�t�����~�ZtK��^�N�4�^(���>Q�d����w�L���n(��Cџ���n�Gӳ#��N)Tp}��L뢜K�`�$��8<P!å��W9:5��5�������cTX���	w?\�������	� F�8��vlBőQY�lݶ&�7|#�G=eE��oQ���Š������w����&�l\=U+��߻3m�����V�[k$�`�+�NLKF����+���3Q�A!\7|��K�/��cj˕8U��b|�]m�(�d�4Bp�쥸L}�T���+{�~�WDpn�Y�û�S"��|����n��#U�8v���&�*�D�8�dm_�Oy����TԬ8r�=�4E୨
��"h���rH�@Z���M�?Ǔ�_I�	����#��	�h�-|������l�������s���N �༎��
�'0~��iloS +UA(3�R+�]���U�[e�ND,o�6h+��5��':IT��#���n��%���@ߪ��6FhdS*5/�b�5}��p�i?���� �[��e�ם�����W�R�#�R�/1�Jq�߮4}U<\.���̳��ꌥ
����L�H��b����<�K.D� �,�M6�����~�x��0lF��λ�y�����Ρ��ӁF��^%�S�+-T��*5���%E7u��Ep��Jy�=:a�C:V�� �.�%�*1]����3ԇ^�c����G��_��a��՚��^�{A��e�K�gv�_��2��(Jn#��ܷ�vƼ&f � ��	�ڭ�OUӑ��G�9�i#t�8�����'Kp 5xj�u�K��e��4�d�Օ���~e֣�#ӛ��2�mz�R��.JK��~�ㄲ2��t�R����;P]�ۛ=���E��p!�A��C:ic��,�X�$�m��� ټ}>n|�A�i��%��I�����OŸ¯�o�>�%��9_�}F��-���\���_�z�E�ިkJ��R��Π��z)������H�N6�)H!���Wb�F�c��0��(?�o��:�7�0AA�оZ,Ȁu�������/y�W���-��c�7�¯�ᬠ���E`��KHr�n�� 5�ų��1��n�c�V��$j^�#���$Ը����e�d�\�//�r����[���&A��?2m�ͅ�k]8Qi��)���G,VF�3���3PL���t���,�o;g��7^� �W:�w�DG?�_:\��Qч1\!�����v�{c?R��������b��~�k5��4��	���0�J�B+�O�j
�{|va8�04Cd��H�;����:N^�Hɇ4�Y(���x�*NCN�d�Hp^����9����͆tO"�!�+���)�%�ή�Ǥ*l]'s)].j����.�f�;n9 �d=!x6�1#�Y6�2b���c�Oe�ed_2Q�i��1���l��.0�����pp������� xV���ÑTl��AӃ���pgC?��:�'�n�.��PU������ɂ���C�Xg�mz��J��#)x9�4��[8��VR���u}�S[efp
`�l��8�+�;�G!9��b��s~���.~��O91N��g���娞�X[O�{g����?���|�s�!/��B�R+�}{��c[fȟ�ן��%�>��l���س��p��=2Ҫ���1�[���N�v4ɼ蹩�s&��3�`H�1�?BD�� ���ئ
S��� �;�<�}2Q��z��R`� ��J��N�� ���upи ֬�C��_#� ��LX�U��E2W="+��ؼAu���}Y�:{*�E�xԤD�%����w���@�8�Tҽ�DoQI���x�>�����h�-2M�R�ܞBA"bѫ>tD}����/3�<���R���a%bn��e�J��_޷�n�����2'�/-<>A�@��!f��{��~�j%�KPfO5����n6|ː[��Z���6�SzX78�I�$~r�v#x�Լ�7s���^�����'���&�&
�Cd�oj���'Уņ�:�.�w�',G.���}��t�>Zտ���\Q��s���吶�����v�`��[�Y�c�� �+�:,�%��<=� �����ZҠ�,��ʊ�Nv���b�_&Xy��:���d\��x�
6���I�5,H?�=�+���r��4ܮ��0־����K*���PCǜ߿��Hz��D�bMp5��~s5SK��̳��I	G��Q����1����� |@�6�8��b�g��h\�{4��e�:�jj�c��|*�1�v��Be�~GM��P�`��#�-��E���	^k�Na+h:�wI�D��՜�qsN�{Ht�a�C��|��Rr��C��P����#��F=T�R�I�S购��B�k$v)lt��>p�p�3��K�E�6s�����Qsxv��I�c_?J�)n�)�7W	��bað���	�k]���������x\��sP|O&���y�8k�����^��L�壘��f�ZQ\EB�o@����|��j�x��
J�~���t����!4ۻ��h2b鶹����)S2�/��q��A&��Et+! v�o:���0Ӧj�;���9���������Tl��������*���~� |(���j��2y��~ t��icFU���>ND�P��K�К�X&��bV?���KŜ�.�s&TUd����"����d�6�H(y*�mtN���Z���]����+����j��fOtqty��E�.���V�d��Qwl�q38`pP�R��J�\���hT>�é��C��f��.���b��~�^�����
��
e��[��Bf��1���O���F��Oc3}Ga��2�:���YH��" ����*�b��%���ED����h�i��,��s]L �h'o���+��c���ڒM��c��*�ݜ�����_b���U�(S�z�,#u
�"�*T*x2d�mң�nn�|p$���[@�6��0�KA�`
�d�us���5�w��[KA���;4 S�g	C�)$�-4�h\�o~��Ϙ������9//T=X�4u���=�M��[	A,Jjg���9���V�-i�whݾ��[��)����XN����6318�-�
��C��JݵCbo���J��Y��[�c��Jw̩�U���O�f�k����0J�0��G����W`�d��^�F� �T�öQAG��%r�WI1MP�:!� �����,�։N���?�����[��ǔG҂^׆���/�^�P�;^;y�´r^�#�9Y��i�tYc@꨽FM!�i�v�׋/���ޔ�������k��R�6U�������|i�%�\���V#��c�T:2���������󰵭��e�7���;�q�"�(�W�Y�LFK ����f��%uJO��=NI�:@)Q�e��L��[Q43��u���x�D������v�\��%htr�|ۣ����SL7	M8KZ�Q��:7$|��_�bw���m*��
�`�dn�D�ĸg�Z�Jj�-+��A4�U�Ҭ)?Q�2nj� ��/{��0�N�v*��2� `�_	�kH�������ጮ�d�K���1�D`!W w�|>?��e���9��+8�cMȽ���$S�!Da�������P��D��碁�fؐ���J���x��٭��K�E=�؋_�`����ֻ*_�`�C%�#r]bG�����j��1d�ܶ�e�A�1DR�O��CH�%��oۍ�%<˿*79�Ʋ
Y�Tu43G��N2�NBi�۬�^7��u���.�pzA�ҁ��m�NL^F;�X���F�T���d��C�@�Eb���^/�S�E�y(��d�g��73�1��.��H���X�ض��F}Q�.����嶱��fb��	t�h�D����TK4��ޢ�SK2��!PQ"I�5+W�;oJ����\����9�7�g_ӡ�)��f�����bu16aM��������o2~Q76��O��):k�`���;�W�O6�w��ȼL-i��A�"T��
��a���^�+��#\�3U�V��m��a�U�̱2�a���V��ŐMd3/����`��avX��j�Z�w��w���n�����c+LS���a�P���9����4�ҵ�,��P:�tB%�^[Mb&\l�بG��OBuh�oY���7l,��b�d��n>�z�Z��,{�ggy�-kc�ctp�u��9=f'����+,�2�W�&��b����� 曐��
{���F`:�͆t�?誏B\n��&aX_p�>��6�E� ^n[�)ʵK�����Ek�4�n�����!]\TS=U�4�Z�
�)\,���O��\���&�I�y��.�sO����(G����Յ�K���=�Ja�,]��I��@���)��S����̌Le�~o°�8�5��	<U�@͞����H"l���<��tT}�jݮ�wB��22p뀡:�\�u>˂4�n�>V2�>��=JT|�(n;	G�I��A�(���c��+x���Y��ظ��ޜv�Ճ�3�daK��h5(�R�ݗ+��=d�s)�5z?ۉ��k7��f�bƳw`������<wˇ���Q�%A�F(�8A=-Q'͏��W�s?� �tƐ�xa_� �?�߳�
�
���jsu�Ԅ��-n=83�-�(=�8[��%L���)�NX��ec�&}�j[&�Z�����3|\��!�6̪E�@b9�D�j��2���c��[�'�苹��6;�H�eB�y�~�7�~��J���/?$�ٗSy�A�z����<Y��z],>��2p��c�G�:������:�Q����;��dD�K�g��FL�\��P������bM���v+�\i�r�������V
��r/�BhXY��E�|j���(�6}�@U�u}ƦЅ���B�^�j�4U�{���oW�^��.&S'��)�����]���xr��'�手|
���(�"�e&�a߶ԧ��z�t�P�Bk�^6���a/��+��j�!J^T� l{����"�7O#�,����8k�Y�w�