XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��f�;:|���z�Prߣ��O.(�#kkJ�f�f�d��F6Ͻ#��M��{�S���K�6P22Wwwn�����O'	]�����,E�\�V9 ��m�:X�x�+&�ѐu�6�`��궝>���6L��˰��LR�֞����x�2}��M�B|o�C>hQ-^}�q�K�kgE,`0B�j`�&�h�3.Y��Kq>\��t7)�9�|Q9��tJ���޾e���>������V�g��*��"�c�#i��r�'А�Wx�y����}��,�7�S�?��ن�E�tM�&%�r�Ș��[l���]Hڏ�ںB�u����/�X�"n-�5m�<{M�.F�.�KX<|UsOo�H���^�B\��;��2g��jH���@S�����>:����P�`�=��w�!�],�=#����cpH=�k(�M�,���l�F��e��B衝̇T���D�"�/�($�F�_^�)������_O��Ų�f?1�%m������(����6�X�2�ZԜ�=���C����9��P�Ł��Cā�?D���A- ��lNʲ×������u\����T���AY��9a�W�l��<�f� �n�@�������9?�PfY=��U�ļj�S���צd��(�5=���!��6�V�wq�)��D�����9rŐ�'Z��;%��=PjV�:!s0�1�Qm��9�hFys
�E�^�n��]z8 �!Z�Z7��"(���si̘Q�[�n���XlxVHYEB    15b2     890��,�o��I�\�����B�<���V��i���X�����ZG[����e-Ǣ�B|�L�&K�(z�G�o�هN�m�C���F��m���u�m��go��Fdzҩ&_����Ȱh���"�NH�!�.�j�����[�1l����0Y��,d�@��A�E��;	{�N.�pz�[��oF�?��ŋrǉ��Ҕ��^q F��!7�!�3�I)�"p��-*-'-;�rń��R���ɞ6V��rɫ�z9ZT��v��X�T��܍� Z��ux����V��:d9��D�9��������c���?��L��dһ�E��[PGt ��R?\��v��Xo�#/"��8h�����F�!�0	R�5F:�D�#�RP�D�.K�
�[�i�����p;��} �`���� k&G�ް��._~~�)�c���Lg��&k&:���7<���F�'U�TVBk���iv��ee�e��w<.ڦ�)aj���ۈ�ƙ��\7��'K�K�K�z�G�lG!J��K�RҰP�۽�Ϡ$�*�L4����d�i�0�k<��2)�������A�J�w$MY�f�/Zj�_�[��\¬F&q��io^|ptT˒}��!!��CT�f�Sp[�&� A~Ĝ���'��71�8lw�����]�b�m�^���wk{��b"4�p� Sa+��x�+�O�쫊}%i�͈]�;1�[���
�{�*�:���Up��X�+/�9�H���e��Z������f����\��ל�/Y�-%��w�}�Honv��d�تkN9ϙ�+�'~��V��{GiD>�����g�xT��>���Ԯy�/�������L���&�����e69^S�:h' �Ky�r;�;�J �Јp����.�{_q��|׆����;ECϞj%�T,�;���14Ԁ�j�h�Q�a.�X�`w�.�L��	Bq8�Ý6S���aYqr��ѵ��i�C 4����5|1�3Q�Du�)*��Q��F���q��6�|�Q��[+!^%�C:�(�)�w;�Uh�ze�#�(�⧾��)��K��_�h.Z�s|�tu�B�J�(��L�$３�c��d7b��1���|�Miu���5ӭ�O���A� ���u�p�;5Քn��ԳǏ��i
%�{�nT�`z�e�VMZ�*2��.�����>��r+�����{N���y-����sD��B��0����./����@�1 �I�9�x��)�̑��8��(ߜ��7��>�)I"������!��✿}���&�~6җЀ�lq7i�]W��l^<]8��Չ�H�$�#��'XL;0�����D��e��n{��&�F��#��ƪN:ף�g\	3w�k	��O�,��lX��zk��H����%��C��3,��:��L�E�{P$���񓘓�a�W!���{�<�����B�h���]7S�?��'t�`��7c�2��@�?��*=s8�|�+�7��+%C��eK-�j7�[.�~�E��"LJ��A{{�vΆ�r�t87�y]j4����O�F��/�w2�k_Ʋ���ki�ʶBڱ�!�h^����ĮڎҢ'HC�Bh/���� vs[�ߛdY�՗�b���%Q�ڃ7���9[G�nnm�K�x�Jht�$�>ynG�[�L�{�(;n/��pE)�	A0<��:�R(��N�h����>���wN��y����0����zȃ��m�&FfT�,��/�����!?�-�Bi�w#�ٍ����2�KN<�&c8V3�|;�'���s�/�͐�?��i֗7	�F��C�6�w��I��L�S�F	�k��V�HC�8��퐄��v0�����NCj�3�g��W"!���~������� %=I�Ã]v�ᆱ}&�1��j��2~�������(B�6.>7�Ĝ��㽆�V@_�
��bi�=~X��9c�b�E8�'(��N&�Q�JG�0����/�ƕ]��`��#R����9��LNڦD�q[J�s˴�n� ��o�����E�\i�Κ�ٴ����*��u�BV��^�+��}���4i����~e'l�sU4�x�e��D�a�,w�c�;Xl���4zw	�} ��oQ���$���K�N����K�