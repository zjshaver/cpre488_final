XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��?�xy&�<���J���y�S���fX b`U�iP���B�u7�\��c0�Y=�@�x�����*���0�1����ח�����a�Ec5�J	<�*\V�1�eo=y�v�'e�]�a�'��&��|*�xϪ!z����p4^Hɔˀl{�1j�y��
�9�)�Gd���ֽ����L*ɐ�DR��z��L6~���݋9-������qv��o��fa�5L��b�>u����W4��ѡ[i�z����OT��[���M��7��
�>a��h�	֮��TK�M�����W���v��*M�~������R�<m���[H=~�oB�~��G�G&���[zϤ�a����D�qp��s��a����}��f �!�&�����!<���ن�=Ú%�%����x2�+���"T���S��/[��B%!%W��X�ȭ������yP�m8-[s��e�/��:�{����Oʸ���T���L�u@eck�p��\~��H��rr� ��ؽ��ju�ֆ[�ʏ�Hڣ�͑ćb���N�U�,����>N���Q�������,%g�����H�����p]\?qki˵{H�-�_����S���P�kA�`�~y�tV��S��6Sn�K�S<�Vl�����K�=J=�R�k1��?��U��eFr�/X�QK�����l r)FOwl��zz�f��Z���)��&Z��|!-����'�R&\�k��ğ�J[�8?�x��.և�+t�0�^�:��hW)XlxVHYEB    290e     af0W�ͨ��xS��t�t5�)�ؽO����	�Z]Y�3�偕~2�ޅ�-�=,��-]���3J�L�0N���|-�{X���|{�_�ˎg���dT��_�I��өWj�!6T����Q��7�H�c#��(P���B����s�����g*Uw:{c�M�L���*�Δ��;*�3����:�=�s�q�G���M�:�'p�H������!���Hl����iA�um��+�P��M�`�u�U�+<>u��t��~��ȥ��H�(vK����q�Vc[A��|B��9]��ݨPrq�-!D] �$��1*���4��wL�,�bH/��d7��c��M y*o6!����b�.-@d:t�j�a�nf�6�}f����i��EzB�i쏅��t��/m������W�\g�08���K��q��8N8���@k(�p*�jj��7.>�����������>q�[t	�|DY-�s��.8����R3"`�NN���u}�E\��j�in�	���IK�bm*�ӗ����K�:
Q�w�:ƴ�m��� wֻv@%
8>!���I:oM�n:���+�1+�L�@����Ȧ���Pok�1ҧ�'�?�.����$�#�h�k�i��L*�YܛёV����0M%>wK���^!��!�7¨�!�b����
rB�آ)�����~��x�EV�Z;�vKzb͘��4�����9�L����_��sZ�n��5��!}F�!"9]B��7��)>���ꉷ�~AB*�R$���Hu��o��s]¥�T���,os��P.����hуmS�ҁ�]'@_��V��tMER��%b�-�C6$��\�)���IJph�sc�sPZH��j�E��5��c�i�+���C1��پ���G�h����<.��@s�(7� �vu}��J�r��!��v@�E���M���+�J�p���� ���я<�F����·��+�g��BsU����^��n�{_u�D����[I��c`u��`S՟K|G��Aj�<��/�-8�A�>v��E]����;�>Lh��S�^�9�E�|!.uk�M!�9���Ɖ�F����� `��%Ihf���"9	���<�I3��ћ�/�`�}i�����訁��&F��U��x")�`�M6:H�w�Q���FK���g^]�9���O�[4^ 9�y�M������F���<�>4�y��C����V�c6M���n~��Z���E����[��qT��i~��mQdQ�sU��k�'��n�o?�C�!g�es�̀���}��)���5|�D�O(| �ކk������e�ü�u� q��W��(G���;U
W�}	�Di	��l���:9��&Qp-J;}ƽu�~�k��m�`�BL� �J$b(Fi�>�<Og9*�Jk��d�N�96�� ��sC���.h ��~�LT�$gԐ��Է��p�����#���2+T�(Ҳ�g����RF)J�,���Ζg8@�J䢋"�ٯ�+o�
�	��q��r����2����cw���zX���t��қ�.���;�X���x�ٯ�њ��z�I���~��)!�Ϝ7q���2�l[n 2�v��H�>�X���E����{�g��'�%,��W�ehi/�>A$��DE�J��ܰ�'ˮ_��z��UH�6}]%��z�N�����|وC~�V���~��p�����8a0�k�9e'��r����Q�9*Hy }?f�ocn�$��S �'v�4�*��RB���el�$���-�!�]�7ɋw	bò2�ӱ���g�w���woM}��
ڵ�q�r<'3�C1��t��2r,yB�v�`��/�+G���q�H��,�����^���U^$�v����_WP��'�LIF�tsostւ$���'�K���V|��a����'���� �ە�&�����F��Ϥ��Lm��LJ��������gt.��	�l��w TOJN��З�g�R��/������#���\#�ݮ+�҆Ml1�ɸ�G�k��	ׄXmg���n٢I����uD�o$�MO�N�3MK杺@�6A(��&! ڨ�3�S�jpn�T�y�n]	C\�j�t��K��>:t�U\��I�~kuo��+�,9{ �7�j���G$�iDcC֥��˼xy��_�^����yʈ�a�{s �E�|�d��ɗ)�Q�h�?�:*�o:��E�w)r��
iM�,n�ax)�f�4���|Z���PnnBPr<	��^O� ���U�ʐ�q�Vkaf����LD��-�ANs���A����&�x�S��ϙl\ƂC3@/|h�ܦ��fl�v��h�q��)�`)����+��!�敕�:�� KPǣ�v?��/P2�wy�`!����B�GXw���|\s�F>-��}���e>�������n���$���@_LP|��
�"I��s�&%K�<�+A�����:���q�s�bt�M����U�
����
�w��K����Ӝ��'2�	� �o3Z���w�t�������5~�'z��Պ�����*!o�q�z�3[@ăuy���*d ��ya���
����W�`��p4�w�|�W� 4q[\��'��Z�A��op�C5ĊM-�2�����!���`�%!�- Y�o�m�#���A�f�DV�{�m����{Z���\3�nP׼���A@ԁ=�'����	{�?m:^A	����.㋏�`��=+`@j8