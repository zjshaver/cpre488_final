XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Q\J)D����H
_H��pµ�*KD�v����d/�eh­&>��Cs�Bmt4\��@'/���s�PA��Ԋd�MvXC_T�`;��.&���]F��w�S;Z�[U޸�ݤ:K��n���=�\��Xsz����*�M�9�+S��aYed+?��2����`I&������Raw��c@L@P�I����Sۻ�1JS
ǥ�#!#(������8�?v<u�s���-s�U��L ��U(Mt+)QeJ�Ę�2R�S�b��.��]t��3��3��h<.N�,#7T����d�R�{����o�M7�s��Z(��q����3��Z�ff�}����d"�?j2��'u���X�)�w�3WGC�+5'?�̡a"�d��۷�!Bj���,a.&&��b�%%��?�������l���J|f�2$tr����߸� �:K�l��x�[�j�l-��ơ0cf*���Z�����j�w��B�K��E��+��)�	n��&�'�6t
�����8��A
O�_�_U� w� ;9�:`��D�!��*P�/� =|�Ur�R����l�(cR;�%g.�m)�����f�^�!���B9�~K|��U�(S���_z��퀍�{M��i�8�2>�g�����f��%Ո��V$b�0m�f&��3UO�*[�F�I�ר��� �oWSE�Zu���'��C��*L070��#���3o�Y�;2.�w�Ϧ��G[t�-#&pQ���W��V�N����`��n�L�ʩ�XlxVHYEB    70a6     b90<B�����v����i��p��KqAi`�71�G:�Ԁ�X%�����=�L8ܐy�k�����[#�KW�1��]l��m��j�IW�o��\�+��K"��5�t�jkǶ����>׼���&,7~� ��o�a;�ف�@ ,'�tn"�m������4jA,�ٯDa^���`�����k��R����0�OL��3�5�l6���܊kpXUß�|o�����U����O�-�*{Mx�+x�w��`:�Jpo�b_�	�>E⦵ߗ������ڇ;����.�>�7���{+Qh�b���5<��N���o'�|>=u0���?S��á`w&�0���ԘX[&$t�il��$�<Q�Kqg�+L���T'F��Z��EQ~����5<WE��IYiP��[,e�ȝ-4"{���9կ`V�::Q���sO������K�v����&�>�<��{c���#
�/1��$$r��[�������v��0Yo����월]Rq�K*.!#/:����ޭZ�KR������*lM׿�ݽ܁5s%�]�D�]��?���4��Ε�~��@���z���ȃV$�g��J�c�ٚ%�?���S>CJ(���^����1����9�s�p��n ��IL�	��:���ul]Xo���C)~E��T�G-�(����z`
C���CCc��_�%x�y�36�oH�4�[��3�	�e|��*&�hs6�D���vҹ"m����Q�N�f��G�!C<,���F����'"���@��v�ܔ����vsY@)ъ�H���
~�
��m�q菎�Rޔ&O�'W��#}�O��P���{-K��s����AW���?1.$��0��D�i�m!SP��UJ0G:�Y�/9|5p���E���u���s��J�wp&�г�
��;�p�Yr��������:w�<Y"�����w��Ӏ���3�k{ON��Y����IhR|�G�	�|�Q�C�&�V�C���/Nv�p�d�6��C�m�����I�D�;?�x�+��|Nn���A~�}.���)4B�5�T�4�v�f:"���s=Mc3�����o�*�?cL�)0Bʏ��v���C������d{�xf��4Ꞵ3���\�@x�$��tD�T��{��c��î~~��h�|�b���A�b?p��eK��0Ų�A�ڦ���p�6s�2
@�.��T���/�*K�4��lCB�"ΘË�V�@��s2�(c��m%`x/��;��C���#�<aF6�	r7R�����RZ�Y,�f��?Õ�I�z�,�4B�4k�Cx��@�i���{����%a`�����Z�n��HE�e't��}�yu���w�:�6�Fwc��ڍ`���:�`DjC�+|���(t�	�X�K�:�Q[�-}R%�2�	f�d+�<�WA�8zi9h�����DL�}�\	� ��<A'AT]�#���	�R;��d�4G)EV>�F��������`�O��<���W��׀�׼�r����1�)�'q[#1W��6�O0-��ذS�̲�Cb�VK?p�Y%C�&���6#K�<��=`�{j��Si
�t�#����:�~��a�E���{�!E����h�u^8�Q�*���t��\H2����!/3��7 �Ft�p�G���r��p���՟� �r+�l_?�tb�P����u�]RX�G��,쉘�Q��w�?4�<=x�!��nU��h�:�帾k=Ҧ��w�OP�lܜ���'���-��_�W�P���/��c"!G������&Jj���O�V�y ���Wj^�\�릠��1��%g=%Q4<�ǒ�r�%L�xv�q����wSy��a�� �
�[�V$g)BP�،�����b��&��q�$2wX���/9MJg�Tmν�S�z�L�Z���$��y��2�9�0�^P���`-�[1�[nR4����Q=�7@ I�M���o��P��m{���&҃!�?R�}��
���`�ϡ�3p�
��7b���r�	$'@N�7q�ʒ_)�dDͪVz� K�
�����
�)�.pf!����!3=�9+IG��]<[k}O��K�o$�#�?�������s[�7�ؤ��\��SJ��X�[��⺺_�Y�|����S�Hn����s��R������̀��NFuF��q��V@�>��M���/��V��������0X#he/�S����^	_,ʪ y{�#��dh�z�h�*�gh�8��<�`j/��+M�!X�ʿ�����惴eR1*��!�ecQ	Y�;�� c.V�w]���1
�tz_M<�vSh�!�B�r� :�D���nm8�y�!RVi�dĭ��~���~+:�M�C��i����k9��k�Cl�(#k�0���_��n;c'zu���C���E���>�(�r,	`�3G432^ۨ�ٝ�N�Qy�%��c��#�{
�5�Nr�6:m��t�}�Ҵt��>�>3H��̬wr{��(C(d��W���C)}˿�03�w1�����a�ڨ�_�Bbļ�f��k3B-��7��BF׬�A�C��O���ω�e�eU��PЈN�v��ސ�+���2��F�~=Y"��[�q����u�x�ƛp'�ʔj�8�HHP钥��_Z�%�m��]�<g���Q�_�H�9_���y@���Ǟ�G;��ޜf����^(����.%��5��!]�G�e��b����K�1H	 d{��p<��l���,ѐ[:��n�f*��!��U+��l^d�ΑzcM�Bi� 9�Bjш����7F�U�Q-G��d�H�;��0�j�e�oO��$)��Ǯ3�� 5������Ӟ�5��}3�"dݫ��"G�]�l��((٦��<L9X�>�$��1g?A'ދDn\a���B8�e'�L�k�G��Jpr5��#�RزCt��Kǋ~3�{��6����