XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��C'���Z���cK1S+\�I^Z���z�Y�E�����	�y�&ҩ���0N]�h%k��EH=�]R���U�E�J�{���ٱ`�@3�ȵ� s�_*�b�}ͳ R������3.� ��p��D.7������wٻN@��4U�9�M72-0� ���) 6#b��Ǳ���є�h��9A=�;��b�??��Hn
]%S��V,����P����c�l"�xȓ~jm����@�7���6�=Dۯ�|��U�嵭�&�g�\��
��O�@��j�{k�JǎV��+7�Q��e�b��{�}P��:{��}fMR�-93���o�	��"n�8���\���q�"@Ty��C��偰�w
�\;t��fd+�-����o�J��ȥBT�5�mh��g"�%Z��g&��S������U S�A56Zeb�?�'��q���x�0y�j�ն���ؑmM�J���<��Klq��Pk$.���l��0֜�U'L�&]�G����{��� ���"O��'��Ȗ�z�C�����M�k	%�O�W���kᜀ�㖂R����qRJ��~�	�����[:G���L_�����X�k��?��cPDX�8᭟j`ȱ����f/ĳy�s��eD�f���+�U�cZu��"�@]��*e*	�]����S���
��/��lǧ���c����l�n�z�c�=�8v酲t��.%���k҃]p�o@D`u+�}@ҩt�¨xFuq}D�U��	���5��K1ۜ�#XlxVHYEB    1a34     990�أ�ڣ�,�X��{c3�Q��]ua7����� �xS���V,���
�*f5p�oEN`���P�t� [�}�I�� �"�GP�J��'�w6cV�g�\�2�~� �$�:��q2�3�| b,�(v�Qp���`�n-k�	MO?y�	�S�����a�d�g{?zMbW75�>|Y���C5R[��Һ�$��T;��{��
J"���&���ci5i�eZ�%i��9��MlQ\Ƽ18gc��	������$</nn�$�<��DT��`�2�o��>6��v��VtH.���6{�e<������Z���`�T)����3~4�E�!������"&�+�!%R�V���"ʒeo�{���}o#<��|tt�/�0��-ac��9�GO�a����ɪP���]ߦ�e��~�1��sA����jڣ��'w�<O
��za���Y�|9ב�0��A,Jq8�������7�P��	�TeS��"�9
"��T�a�b{е ;��EP`򋳤I���7���$�>�B�p��$��ǀ�(%�}J��7�4;2�`y�H�Q�<z
���|��>��5<��D7-ю�L�Ӯo�B^W>@�_����	�e��Fe?
D}W�/`~��t>�iv���NT	�3�T��	(1�`�Y]��]�sV-CΏn�gw��铖/�R���$U��9�J�RR�?����`����̀#[�2aJ����)߆����,��ұ��ꛀ׎G���{�|﬊UԲ�-�8�-�kms����|޳Oĥ���	�Y]�]���P�`��t�(�R+���JX���tAL
��>�C> �N�b��6�p��-j�:SKX��ʶ�����"-4Ň�˥�i�?��0�u׈��q���h�|�[�U��!2���4�܎���W�2)��si�-*���dS�h�gɆ��ƹ���o~"�"�,"�R��{��T��2l��d�H͖�ˬ@B�������L	^�Hb��w�ڵ�7d����+��)��(�/�?K�i2J�aI9Fcn>�ŀ��k�~��SY]X11�����$�Q��/����
��Na�"����,ǃƍ�Kwh�<��!�ׅ+c�=���f��޽(y0�8mdCT�b�g�������}�P�K?i_8ِ
�a%I����ệ�b'�?P����q}�Z�o���jg������抯�[�vKʙ4³ ��������Y	׶�j$	�G)�Њ&�����չ��\�R)
'����(��mؘI��ofl�P$������s�C�EPѨk@:e���C1�&U�����{v�3��qD�3�T�E��9E�{gW���l���o��Y/B�������e����{���%;��r� U���?�jjy�.0
U�Dlg�%}j� Ʊ'�F�
ҫ�V��}w]�	5HdD� B;$&e���?�������~^��c1}WW�2���Z�ߪ���[�YQ����&r��;�ݢ��>��i]H��a�P�Tǎ"�%�Թ��0g��*6�c(����|�#���jN��f%�}x��K�%�L�-�����JNr��g\AKl�h�C�7��I�������d?<����nl�#��6��5�T�+� �y���vܘ=K֧@����
>��n���	Y�L���gP����l��2b䒀Y��.����a��;���_�|�����1gA�%�՗�
V����N����w�Z��n�UZZ�^,�kӈ�Qq!��/>x�4���#o6�#����)z������#�S�dG�7r�l��[�iꕽً�2k�^���/�.v�"c.5`[jM�ѫxd<W��A���B}Fn�?fH��W�5�؍(�y�>�]�lxU�F�ڰ0)i+��O�"�q�cP��f���0�v��������t���Qd�q3�'�g����PG)Z�.����p���2�ꚃ�� �L)���m�+�8�甀!� ����]��f2aۭv�Qk��8�}��ljh&FgE،o-V!�G4>�h�6��V]�mOC�Xղ�	H��Y�����-��:�d@X���W���व׵�U��C�ɚ���{z�V��̍آ7� &�{J�1t��^W\�p�Cl���g�j'\&L^ GD��h� �+� h��Q�?-J]�#sD����4��(�D�X �"��O��q����o���1�9[�5�w����ĕ����`��j
ϩM: f��kn��b������+�g�1��xt���o�l�A�-��T&*�����4D�dѯ�5�[�rM�k��0�J �'8��39sL9�JC�z���w�e��a.����z�������g�6��R/��ǹ��۬ce�Aǀ�pv��>�K^�J���Z��1