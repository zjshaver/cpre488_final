XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���}��xp�!��{�z���٦��k��vٰة�������ǰ�J�v_�#+��o��-���m�}A�Xs�U���o�+T���C�u��ODGl��|�8��L+5A�66��>7���,8=��,F$�+WԿ�f���t�Ͳ}Yo�5.eA��1��"z7#�E�Ņ���#  �Na�~˰tt�\��8�,+eK*�ַ�TE����T��a����H���ݔp��5	*K�eTt`\�W�~V" ���ƴ�r���TߍF�&�'���\�����'�!��vkt8Z��BTd��q S�+�����54��I���c����8[�]~�L�=���]����]	�Y[MΕ��KH��"����"��g*jᱞR����v[h׀p��<UJ�)o�%�-	f�I��wT�2�Ee������G��n�~n9�wy2u�y?���4��ٛ��z+�h�a~Ӿ���؛	��k6+%"yоp�rE�ȝ.{�;4����EB5�э��*���UR���hR	�jP��¹	�K7����+$�po�U���1�'ڣ��}D��Q=�@����f3
�1�Z#d~4����'��/�X��q���u37҈m=���d.�Z�g<Lř���b��0J,y�X?����f&>�x{�?hX2y(�_v�:��pԐKK\h�Tܩ��ݿSs'2x�^����K�_~GT�k�뤘���;��;�r��6���������mo����Г}�N��dF�Dws� ΀XlxVHYEB    82c3    1970�N3�>O`�-'X���slo����-2�5w�2k��;�59�W�B9N�CԬo���d�Q9��K� ���z&͔_�Mm�6�P�$�a�Hm���=�N���"FY�nlm��Phh���?���y���%�۶R튭g��p~�r��5嵚/��4ȱ��*����B��B�j�_�_��Z��j����i���9s���>|F���S=����@Ԟs
���g�q��n���!�/�e.Uv3"��}��.�4��������u��C�v�|�ڔ%��rƿ^�n>�l��Cn��Vỳ[�5C�O�>((��y]��(Q)�y����n���	W���(�#U����J�C� �;%P'a8��J�}��*ݰds����������	��u��A��BTh�QXO��幖*�R�^I�R-"��BHlw�0y��'���!��$�D6=�L��-����W׷dḞl��h�Z�9ր�ّJ.�����9O�[~�`b��f�V?WC�R���N7U� ٢��"5���!�}Yg�k�-��}��2UE롅J	Ax:�"4J;6�X��7{���J�#�=�k�z/�Z�ζ�_�D�U>��ű���������=
Kvu�P�����$��;O���ᓰ��߂����1r�${�I���@S��4�\
h)<��G"�"�^�7'l�����%��ThA2��&PO"{cK,��%޿�͕d�3Ρ�x�%�1RW�Jw�]ȸɛ
�%a��Y��z��T�8�𔦔�_"�"�\c�G�m0�e���Y��IH~��<Gk���l-S�ܷ��d[%⺬G4O����+f���<�����
aR�/���5v��B[��J����=���0�^Q�;�Ɔ�����Ӻ��U
F��;�#嗑8F|��5�k)sgl\�A^��J.����ԍ��xq���A�.���?�����fX�R%���{��?ͤQ�8�i�����bX�r�b� K�e���S(6�b`�Ն���=�{���38��rN�WZE�4c�6��Ǚ
2��0I�q}�ͼ�T��ӿ=��qB�dDam�����8�[�Nʻu>��ш\h��o�q����U����i���kή�1 ?;)�����ؘ�p�僦E���ŗ��-7
{p2;�sчW.5���Q�f6�B����ٳɇ��l-Y����a�N�������	�SE�-��u��'_�v�duʵ�e�_l�=f�2 �
���,`%�9/��Ͼ��!������~��) b����b0�����9�fV�V�X'��8�gÙ��fv!�5;O�<s6 k94�@b�L����V��|e�z	��w�*A��Ѻ�:��eP�����͞]O��������Qjkb#�|�va��*:�Z� �d�>�b5J[�ꇼ#G�}gW9}(O�b���u���E��G�BF|��2(w���ԹZ6z��[�� � -�'מ@�;M�c>�V�2&�Κ 9I��T<�0N��������5ڋ���h�$��/c� �=&��nS���Qr�"!�4"���N�7�N�]F��}㶉��� ���i���N&jf��6�.^٤ۍC�u��̵t�
 7��a�?���6�F�� d����,��HQSn�����̀�q�;	(�h��`WL38(��a����� X�MdSަ��g��O������{/����>BZ �QX�f�60Hd����PUKfb68�k�=̋��<�a3c�g���لc������8��;P"�PR�#>� %��U���G��������=�2\�-"�QG<��{@魤�컬0^�f�L�h�+����IB&�]P�K W�m�#_Xo�f<����Ƶ�oɲC,ʕ��~-&ʘףmU��v��]���X�\�ɫ���xLj>�K�q�
:z�L��YC�<^�U.o�``�H��,�ꄊy8O��Rg^X��ɠ�ȴ��32��}d۾?PO����5m��Y3�������"Rs:`���yzpø;n��(�D��.H��j�9�q�3������?�+�x�m�Z�W?�dM�PƂ%zx�R�#�<�Ѭ���c�v��s�\\��9�5��	�����,If� ��=�+�N��U6�\]��o����D��bM> i���i�e�v�8LPo���&��EŶ����77�B��u5R:�F�3�F�Hj�p,�ޗi}K�DE�5�9j��,�Ӥ�~�
������J��ϵ��b�L"���FTYbE�x$��q�������W@n���-JW���	Ƹ}�d*3(�$���;�*G'���;��^�N=,5f	�A@��yR��@�b._�b7& ߑ�X�0T�鈾a��n�Ic%+�.���t�Os�I.k�o\[{Y§�tQ�a=�t���I��N!�r7��`h�a�хsC����l��Z�ᢏ�Ǉ}�\K$�hm^�j�"���UV[��v��^i|�W��7(�ۭd�ڊ�UBz�ç����1r޻ǎ�hTA���;�6i�?�{�l;�R,o�����s[`�ƜƢ���Ǻ�y�l2Fr�c#��h�Eδ�}���9��\j��W�����b��X ���׉e�I^��O�'K� ?�<)j*n�	�Ƈ���l§:	1Vn�9�O �ղBjf��K����Zh���z�1��M̵۰�WNVf����&lEϧn���"�~��$��2��O,(���uwI(g�Hwa��ˆQ�6�� g,����jן�����~K�r�Dʃ���d���G5E����݁	3k���*��eq�W���E����;��u��.����v	ʞ���'6�BD��jۗ�B'��9��Qh�jJ@�h�����x�jB�Ś�Xl��C0l@m��6��r���"����V�i�W�0��̌�������X�j����2	�ւƵ38w�������&I�nb��Й��Ѭۭ���i�Ȳ�\^&����*��%�{|x4o⃀{����T̞��F��k�4Վ����\��C8":	,�)��u竂����AS�z$�6_\��]{a1=�P�}�el��ʄ�� I�"�!�[��)���Fd�M�B8�7�[��L�C�5e �O��˕�Z2�i�6�/����ĎX/CF1�T�y��A ��	�Ļ������K�fJug%d�3�]c0>�|?��Ѯ@f��_�@0�&%"l4ח��O�`�h"(��cD���h��Ƀ$
�cs������ڌ�@�ЇXf;x����r{���_�).�򶦬v������e�C�l\���8Ă�}�������k�8�Z�k���"��9i����Ǫ��t)(*�e��{�_�� �d�.���t`��)@������n;�R�5N4-����Lq3hv������Cɥ���U�H����MY柴��%؋�W�hH˙�����A�:�16i�Z���B�[^�C�@^�l[�cUJ@X���A��4�J��V1��n�ip}��a�)X6_�g��sy3%��\袜���VӰ��/���f�sQ��vm��<8�g6z[#��9e� �-�󄉯�[#n��%�yv�.��������.�d�D�H��['��vq+��O�<Q�[��8�������@�����>��,�Z�ҰE�0�m��H���ӛ(bE�����u���$22
���)��;GK��K����J�XI����q�����р"��d�硌�����[`WsA#����aF��Ew7�!Hp�s�c(R�m�4�W��t=���3ŗ��Ύg�
���*:|_-��D��'$c���;���
��@P���*���;�p�I#x�1X*o��A`/י��x��nX�4�w��u�끠��'��	��HG��M5���S���'��5�.ܵK�?�M�5ķa��!J�p;�Λ3�=]�d�rH�""���u9l��j:W��h9׋��[������0�)��6�i�cg{������6���Nx�c��_z�5렅s	2y8��|��n�s�7^5����ș���y�*uk��~�s�01FV�y~���hm+X��&+@e���*�-�;�nW����B��c�Ox�eV�;ɦa[������s��
�T>�3U���� +���.��2���G�x��S�wxy[�0���L'�ɀ�)^�����y���j랧�P�m�?�c@�2��do�(��V�w�RF�f~}�2~���F�s���H�� sW�A'J]L��X�Pn�M������q���A��JV+M]{��[��/��~���R�:�m�S@� �~���O�ê�ɹ&9�)��2A5�1�wCWU���U�6��N��~(D�"�h��Z��5?�Z�w�{.��x�ڃ�B����'�QX�y��1��5+_>��L(8z��������a�x c����c��E���mk���DL��,m�֖�.�E3��?�=`��6���� :��ê��G��>7��f��m�DoMû>Pk��A͍,�26G��`�a�UABRB����,̨�OHW�Y^#oK�uȠ��ӎ��<\�7��b0�M�pIX����3�I�� #yEZwY��q�w&��f��ِ�7b� ��&��/�
�wc�fػ�s�S��u���o��Ф؋���;�yK���## 8}CXWҺyD(��t�Lg���G��|�����kGW�_��[���}$�*�򓿃����|mD�Z�|�7\i>�z�0ͷ_o��觴n�Ih�A�Z�Z\L�!Ƿ6��6o6V�aY�ȿ�\x��mK٤"�Q�:��@=�kcO*8���\� �F�rO����V�j��fKGJ�j2���w�8aT������ϝa���.�5���.����ꅭ��Վ+Ȭ���f��xm)\���d�]���#��R�9�<�F$NzK{t.� �aܹ���u��X_r��B��'#�~�T�vwo��d`,�Uc�)���0PIg<g�
�n��$���`����pA�pa�q��lW���Rę�7� ��c�bU�/�U�c��f~kxN�%I7�%t%�������3�Aa�����l�5'��ĭ@P6|LRL��*�Ԉ�0�_,�7(��kd�C6����(5��A1�E�-"�v���������ef(0��z��;E�ϸR9J�Z�u��G��XՑM�d2E�:E史|�*';�ßT�<{ ]��믔S �TZ��B�D��X�*ISZ�!a� �AL�/@��A��ǉQY�wT���,K���X�se���ס�Џ�b��Ί�J{�t�#�]͐����ọ���g��(�r:
a�T�a�
>ү�p?@�_F��<^�@b?��߱Ev�]�7ř�����Aݏ�c��3V!҉V����U�V�����G�z�l�G���m��
�����n���-1�CR�`�������@"�������p!Z�����+p�m]�"U����ۢ(L�F��5�����\~�
��8[ ��&y2?#/I�E���4����Z6��^{?��D���.����ߓ
���?�a`��4��Ma�E�Ї1�c��S��Y�{ɓB��9$,[��6�D�UO�p�Z�π`���k�doW[<���ЈXe�H�Wi�,�@'Ǧ�C]��j�$�I��إ�kH�p�,ls����9
5�Y�$F��O��x��]�w�^� \��p?��B��딤�qJg��t��T���mj��<�,q�����C"q�	[�&ne4�u�KX���dĎC�wI�%�����} )qg:A9B�3'(� =Jk�W��яr��N^��aqԩҷ�x�h6�F���J�����u��8���v˲��E���̼Ds�I8\�IWO�UoyYN���+�F��$f|�(X��/�I~]�s���)�)�gߍ��k�eo�}`�2�)�`ۃR�0��AJ|�_����f�P�A��NLP)���T i���`x�ρD�'�
u��)A�ǖC:n�-mѺ}�G�hR^��H��R�����G�
���4��DS|5�b����EC��p,>y$�P��u�ߡ�Z��_j�����ß|m�BKo�Ŋ�0n��v�A����JHe�n�\��2����_���[��N���s���g(O�4�o�U��>��ی���F5DR	a�]�� �k
�z�U�����]������q�>�o� ˷���ś�Ư� ]
�؄۵-��D�x<�@5%�c�h�`Ȣ��E��� �)F���{�Q�0.�l	�$�;�X�0I{]�����6�ep2�d�=������4�_� i͡1��A�7���FDz�����?��>]�ù�G�0%�o