XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���a�m�рc�m�y�c���r�=�nX��}l�Zx����>!2{ئ�n/㧑�^���,��y�kѲk�"��'��*�k<�s���>p;�� ��EH�׻��~�ا6���\��7�.�z�^��EP��P�;ml�-F�����-� �aĪ�*HeۜĄ8�Wv�V�|���LZC���q�	��)o�>��6����:Z��\/d=4-�x��+�"&r�%Mu�}�a�;�ޞ���~�F-�4�^�j?�K�����Ə��$��o��pj�Y�����iQ[�C�BL+{g6E`�9�j'�סy�1��7���:9#��=����uO�o/��\(�ܒ����	�k՟�cf��\%�WJ�.�.*xUNM�
�윀��-Br߄bN�}��S������;D�;ǂ��l� ��	�$�+���'���卶�X;동LGU���6q�uy1m��t��cl�r����6���a4mN�;�za�B�x��lZ��k�o�|>�]X0!U�9v�Wc��O��Y�(�X����-��t���/3e�HeH0�>������e��-�<�:��I��3p��\aCsGجs�O�쭠yd6O�o���۟�O����� v��t!a����֮�&���g��y�����49F��GXW���i)�n�>2b��*�z�=����p-�4^�5�,H#��%�����a��e7왁��2�a tnr�����j�%�:�}��q�A@C ,8�9�-z�j�5�k�:�XlxVHYEB    925c    1a60=��)�r%��4��)�-�������W	X��6�;F�8�)�P�K���i���pR�(��q�y�X��45��U2�Z��lǧ��x�s:�?�h���O(�\��
��\\m!eg��E*TGQ#���+�gV��a��^��k�?�{���r�������F�9���ŧjP�sRf*�aK�8�Ye���t� Wz����f%f���#��n����C�y=���6�/u}��I���&��EZ�q�!t=C��Xт�H��H9�B>�7D�����^�3Z�L��6R�{3[]��Fw
��w�� ��c��x5�2x�X�S��@ƺ:3�B���i.*����;��mF�oO<�O����fY�1�k������
�����R�h'؊b��8DE��΁ߔ-�B��/"�~��s��(#m��a���p��#�!9u�^��>�0��q�����W~�S2*Q'׃��Od��{m���;]����((�P֍tƃ��o�&#�)UZ�_��Y���p�n+@+�&B{#�u����1ח��d��xH��
w��J�_�9AG �OW8�	U���M�LZ.��ƣd��6��!]s�|�m��.Ɠf���g���0�I)�g�U���x�/I�-,WƇr�BK��M$�"P�h�L�u��a�xA���x�{��Q]t	�RS��; ����Y�`��h����W�q�4����{쯖��/0�oԧUY�ҥ�*�~qF�?5r��4��?!ݭx!�^�m�b_��K��^���Rޘ� `+>������@7ɷx[)��"�Q��8�ng��Ŝ���6.V�ıeo��!�|t�h�Α�� 9 �A��	@�/��Q���jW20��ZA*9���\Q�``fɲ�o
2K��cX��_8��}B�Img-�dX�{�E	<Ϻ��51qϴd(tuxI��lK�H�Z#�h�qu
�nK� .����ހ:&-1����'�~� �?x�C,�H��*�0$����;���6���-��8�}Z���ʀ+�@�PT3�`�Y89>����f��� �I�9L��W.�Xj<���d���r�ޓ�a^w�Y��f�%?^��C)��֠0i�V�{TV �~�_�9P��eE�}�`��|���3�A�#�u�����͆�]��LJD�Y0��g<�Я�����ls�*m��nX���<
Ӄ͌�35�\r���
l�C�Jb֞�BL �+��xQ(_�:���u-
�?�|,tS6�	���[�Wn'w<�	����f����~J,��C��̢0��Ǽ���ۓE����i{�"֒�L>M�4��D��޽,J��Z���?��*yh����jLvko2[��AJ����f�N��*�c瀹��&x�7i�3|�����HE ���p.�iڢ�算<��M0�����Xp!AM'��A3_Ce9+`Oz�}�&�����U����U+���jͣG[ҋ�ҝ��-��?Zv
���?��{�n�DY�& �.SJ#Q )6mP������{��GGr��@�+�[+���:�p�ؽqܱrR��Ύ�?,�_eU�Y����u��#%�m�b��:>�d��AcfCLH�:y�Fԋb�M�r/~�X��-���=ީ*j"�*�Eu�\���m�f����5ɸ$�� �h��d`N��2�O�
c�h'��q���N훹	>Ա�y91b�军=�p����"���A00-&��x��Zx��Vˈq �K)-�BI˦���N͝�-�;�{Ot΄�ds�X47�+���S)�P=V������z�Tp�#����(��T�}~�E�PI�WpW��՝Ժ+g5B��ZL�j�"T��x�>���,F��M/�dYj�u �+�oGRÅi浖�9٫@�	��/���L'E��9vM�Y�[ǺC'TN/���lB�C�ձ.$�b���<��r���XǙ��_�V���J�z�F��.w=�cb�-�7+��r��ʜ#�x�N��Ec��z8HBlCWk�Me��NCxk7��q�Ů�Yle%ƹ��'�~6*kM��eI��!~�k}[т6�3�#���p�J����
��G�Փ�e��nhD�N�	0t$�'�_bu�=�D6yK\�\0�E*rB�	�ƾ�4Ą�	��B�ڱy-�%���	al��l=C��\��'S���4[;��H�\����`K��b�i>S5k�Xy�R�9���Ƃݸn�9#��C�7$U�f7��.V�e��H���3J�ǖ^�3�ȥ���ʲ�kI��CO�+�Y�jh����(����|E�㏭Ӂ�|������ސ�"��B����I����ծGW8�~K�;tjn�|p�[�X��9�@�T��bM#DZ����`�G�T��~�Sm8��.E���s��yk+���U=�l�%C�*��e$nV�!�����i�:CI,�k�'��[�tI_�Z���]8�hf��X������p��`	4nt�9q1�i��I`�3�*љf�l���c�8�\c-�� �8yyP����2g�[���J)�u��O��F���o0�[���#���Tm+Pf��O�ٺ�����Te��τ֘ ��i}�/�i���	B�-;�okHQ�MȀ�Z��6�Ht-�&Lq�(Ix�k׽��~W��"��` ��P��z������(fl�ί�'�p�&ݧ�iԢdm�@�T��	�����#�<���}�@ǜ`�k��Psҋc�K	�k���T�_�z��U|�IG
�lu�:W���E�L*�����:�Z,���xh��&�P�#���[�
��"���
��4Lz ��
E�i��ӳ֤>���.�ʸ��#��deFO��}svI�u� nf�9s����u(�v|t���H�؉�]�����I��K0Y�/j�u�ՅP3^Cb�k&�!y�v�RO��w$�2��X��o����0t�k��V�̧"����͐���dQ�e�QX�B����-7�􁱏�.�^/���D�߸y�U����;9�4=$�'i�w0�SO��bZfIs焧0�a��̢�%yq<�*'�2]*ɺ�`�G�z��ju�J�;�G g�G0���`�rO$5��"����|5G�t`</&��kxx�~�tR�bÆ;��;:�U��U�)@oF�5�(1��n��K�=f�؞�G+p��V�����X]���a�^2���Pʂ�Ц~uq���mԣ��Y�����{�:bE��bL�H�R����"o�J�1�ds���&���,���̺pX����-�Q�n���U٨
3wU��x@�b\M�	 �Ƽ&7���&�ۂoV7�YԆ#gS���'�~�ХJҸCtO�)[��
C�{�T�y�(l�!�yL�6�r�x�;2^�vI���)��*�&�L�	.�7��2ޯ��z`��zC�QT0���տP�:n�S[w O=+�sNfӿ�A�ѤF�]�����K'"c��Ѫ�r��5=���2.(x�wۡ)zH���q堃k��L�s)��m�W[��@}҆"2Ƅ%~�<�p�޹�b#�w&u�D��Q�o�	v�9v�x��r�/Ȉ��yi��ޞ��x���XV���srv�갭�<�#�B{ji0�S�qa�w���@���bh�S5�w�Џ��cq������B��C�*���?������BC�6
`������@g =��9����o�d��?�l�('n'(���
����v���&�c{m����o�L���b�Y��Q��lS<�k2�a!ͰR���/#��m�����x��[��������
ȯ��i�2j ���pY���w�2��B��B�%�k�G���ڰ�f��d��R������gg4{� �_� Lz1@aX����)��[�����9_�̜���*�q����'kD��Zb1H!WO�쿟�<��x&�r�J=���w��Ĭՠ[:�.�[��7CO��X�#��`P콮�d�7O�[�F��2���2�������9�eJ{Ֆܓ�H9��MC9�EI�Wi�6)�iYE�7F�8�m�M�7��%j��7/�ސQ��j�<V͟��(�8/�%v6Q�+����Q')	��.��Z?�K�kd ̀�a��	��f��+�&�g~:MR����f����d�0}d�\#�v�HX��>�Z[�$M aN�'���be��"���qeu�h��PT,󮍇T�VցY�;_��Z�+�0M�����>y�4�&���Y[zR��ާ�k�Y��0ۯ.�z������Zѕ�Us>�Q�Y���{��������L�(�AG\� ����U_$jQ?	���T��Y��v8���G���dC�=���C
F��){:��\ӿ���y��u(��0�IeBW�!��=:��
NV¹�!	@f��$)$�M~;�����&��fO���I��yC	���1	�yQ�)�$�;4����nV�����l��[F׀4*�pD����M}��a���S�2�C*_�*�A�{ܘ+�0����@Ds͔v 0�b�dGaS��>]��E��u$������S{6��%���q$Y�h"+>
��C�'�n�ſVl4ڧ�,��J%�΍z@aQ�a�-U`�Nu��PQco��q��K(��`�!�e�8��v��c��4-$S/�b㲫O��	��*����v�y1|Y�~#Bxsl�q���i ���n��GwuI�'��
��Aޔ����첖�R�zmdOfA<7v�K��tWٗ���8��CD1��׫4��l�`;����`z�8�G�2^�6߸�9^h�D�̙��m��E�6]�g(�Lz��I�*��A�U	���,��5�m����u�=������-�6�W1�v~�cO5o�A(5�}���
�K��v��m��J�S�Я��L�p&�����uC��&nN�ڽ��!�����y����H�:��ӯ	����aT4�nਊQ�a0��,�A����ǯaX�"�jU�^��P(k�#�$d�e,��a����k�I����OBDņ��o��S2=x�W3n�?$�
r"x�pHMvN���~`��c8���d?!�&l]̼|	�G6ք���-�Zm���ɳ��=�3��EU��*C�b�� fmB�	�A�]�̀I����x�C9����K ��`"\1�1}�[,��K���:I11�+b�:��!\~:��z���E��Ь�q�u��Uގ���BW;��Ļ��2Mdy��!��m�QzJs��� �7����׳�x�I��j�HJRh
���(9�R��\r���ԏYd��	b*J�K2��i�5h�@��%$~t��Á�M��XN�5[������I��^�[�T�.�k)��
�V=�?��V��W��kr.���Oy�AǍ}�hU豋ܻ��,�
�c����]�H/�.X}����}�H���"��q��l�ۯ������
��=Vٻ���}�!����i.�T���Ϙ-f�^^�d��&AP5&iC��Z-�o���L�cDLK�}�j(<qt�|H"�X�ֲכ���my�6�k9-q�` X�mdz���U��:���Еr!6�_�R�~�h�06(���nk���N���Q����qY\ڷ#w��P��ˏ�%�ݲ��~ޙcɡ�����z��<e���ZK�Г����h�g3֚��������]$?8k��I��:H_�P	%�3Ok6��C���D���� $�7u>y��(�{|�f���hÄ&������y����k�he`
��6��Y�LX/6�Z��f�v��-T�`��K�@TO����r��]�>s���yH���_b�e��W��o(Aie��?�0�kX�&��g`[5g����@��w�ʯ>�����y��I'cܹ��\�Ǚj
B��.�/������������a.bFv�N	`��JY�]3��s>�{��0�b�]b6�1"9,��f}�QGHKL Ѷ�_:�i܍o|/"��AZ�%V�\���%�ף�C���h���+�Oۋod��~_�~�<����>o�������L��Úd�2��g�Nf�����#�g���B��7� ���C�3®m�рE��Α���*�D/�͇`x�WQ)�@0�;����ĳr�1��ۢvD�ͽ<�D��9n���^\�u����t?7n�&j=i��h6�?���T���}����jgB&��#�i,��׬��M�@J9�E>��ʺ��0���%\!ԛ��,��7�9�L|̜��rΒi�#�����X��4�A�04ݞ3�z��-�D1�uGm#pM�:S�B��5bͩ�9� �|qGA'"fƝ~��{�73g�!/g�2�=���=�� X!�Lq��U�ǯ����\V����ಝd�z��˩��Ǟ�5߸�n�1��O����fM��9 �'�a���|�<`��V~�r=��T�ZV��A����cv�>���M�����Πdzps�1��o�ps��2cY|�{��L"�.`uh�ܾ)�/5� �P$�4��v��/ٌ���n�hh�����t�����`���j���I�Ϩ�bt��r�[W��e>(�����)����
�z��h��+�'M��Ձ��ir�δ���q�s�	=�еq��� J]]E���dA���fuo�B�+c��