XlxV64EB    fa00    2a40�N���8���A��0�����GA^�J�д�+6y���sdV�]K3%���sX>�L�D��/rdX4x<x�!Z�H��9Bb��;����5{L7r������o4rl�+"e��ınڂFIJl�"�5����6m��X\�d�]+z7��R�׺�����"_�S��%��K.�Ç�j'�Hj/KT���,��d��+7i���p7��zk���G\��4VL5� �;��0��Չ)�(;O��m�,�9.�6RO�]�w߫Uo�Rb������������X2~��q82!ܯ���_��L���_>���\�:Г�>�l%?�<�A����I�I��������"�z���h� �h��c[ih΃?�KN3�W{T��ܱ:|�����8��Y���Uz9���mD Q&�=)EU�I'�D�;w�.𮢪!NDa"��_�����?g�Z�W+LȘ�!C��V\�W:�<�x��8����r$>$�t��@�J�a��83���\.�A0� !x��9��Yϯ�G�0w�e��z�mL�h$������9�Z��A���fWw�afK#h�8h�k6?�
���ݰM?����/�\�hv��;��[>E%�;`�5�@DbN�Ž�mp#�2�TA)V��[�rjR
%U����V�D[�q��)�Lջ�,�n8I�`
m��P��FG���<�����92SR�X��������-~�[DS�ٖn��pqj8M#O�%��	P~�?0	I6�'����U��e��-�;�<+��F�͵��v��� 2ձ�2�۾���1!G�A��~uN6��y��FvV���uzV�۲`biR��M굽A;w������O��a??A2������'�R^��)�2��_��/y�:��Ek�yԐ�����ptԧ�=J^�R�4�9VX�%�Eh�Ew���A���0�XP]��]k)րK��T��?�^�E��F�Ԩ�Y�ڗzc�UԻ�*�}ތ����K�<��NE�%�iX�d�<��M�2�G�5��^�}R�U���p�K���y�h����!�Ra;��0��P#�fAJy�!�[���.�@6j��rf�)��/�z�<F|ԇ�8���D����a�GC�a���6�J�mժ����<3E{����R�m!5��1��	���2b>�6Ve�U\R_��z��	.$w+�!��������3\��_ࢬ��jb�������@��O�,_��38�E����vq�ѱ�\���^Y�=~���Ѯ�>��kc~Oii�2��+�s2�������� �>x=�	]�&D���d�7q`B���ǋ����4�nj�aD֌XL}H���#ŏ���h���Ə�{�E>�8�a���lP�Oc��!)����Ӕ�#bh��7$T\��+rF���--��HQ����l�ZAq���c��ͨF�A-���$ݢ�t>vt�!=�� ?��E�� Pp�����5�����C��w�>�e*	�g���u��f�G��J_�X���:ȓ�C�T�����P�gHp4rOϖd����o|�3���C4����܍�#C�NH:YD_0O�-;�f���a�9��yL&��#��BH��,�+�`�m��{���;�̶4�*dM�T�)��׏`;��a�_c:��z-#�<�h��Eߖ��E#�/e�f��]@���eDe��v?�������p1VQKR�$���%c�ٌ	&n�\���؁�sI��#�d�C��I��s<|�i'������$F���������*�P�Okj�A���Z�#�J^��k˩{j��ypEK�<�h���ub�e"Pù�D���/����ٰ�
[����yy�=��'ݎ8�u�#a�I[1��*�OH��G�lo�3��d�Zz�c�ྮuu�9uw�[T�_���!��Z1�ѝ$�@�°'�)��	��h�M#04W��h��ig<�e��
k�*u?��0���Q��j����"���^��}݈4b$`e�3�u�r(�(?<\6l�/P�Օ�=F�#��b�tt��ι Yn-xw�ۙ2t*Ǯ�1�o�̱�Y."*��/���OPa��]*L@��e��h��O
�|��m����mfF�>�l�C�2x�Cf���cT&w�gv��z�����c��r���u����yV��VNZ&�xC6!9�5� ϱ�`hAF��Ų��*���|v?�XѼ=���v��=��y�7H$��p6��[�cC���n�p�i��6Vy"���Qo����5�]/�hS+q^v�$��a@����^���u���qgwa���@�&����Z=;��>_��XS�� L�
b�/=;�\]ේ��j,�3��� �"� ¥2��V�y�C�id�����Di��ĵ�4	ZN�=�^4dPP]�-�*�8tc6w+B�8$#E��0���oe�y���6B^����0e~� Is�^b�K��Q�Xt�*ʘX2��XJ] �� -ل���e�Σt�rX����v����Y�+���p�t6?�������`�y�����}�K�3+@6	lD�h=E�����9t3B�/�\��O����ݏ�wD�i��	��J�Te�L��Ao>�h�^�ƔN���1��n����{#���� �lL��N�e�\��^��瑼�j�C̼���0�Ԉf��jE��dLe�*����# �oXpk���@�^d�8e�j�ׯ�_Ý����h��'%ף� F�i|��/.�6�9���o�ut �3b4]?����~\S�nBB�d��� 6zc����k;�gP��`��07�ϔ�?����{FEps�Z�����{�鿝�,%�m�mӿь�ߏ�dY=b�u-\�$�j����#f�vb��JD�+�R@��g����d�|���_��:Qֽm�P7�@m	S�����٪G��j���A�����i�+o���8�g'��y[d�_��j���ʀ�iRv�VB��ڿ�����[!����k7���*d\�� ��&�mh�8;�s��^�~���|S;�2��[�?�޻��UA�"|Ͽ;Bh�\I
��Z�����as�A�R&�����ޓ7U��-�&���J��3���&�O�vZ��G�q��S��hR���zr� � #`o��`w/�ѣ��8����x�Ga(�F�X_i���_��%p���'�q���U�0�)#"�oS�Jo�p���ŵmܣ䷪�vR�xQ �x]zX�|+Ϫ����%ThP~J(�f%y����o�BgS��B���g��V�5���bL#���`�{$�5�!dґ�Q�$Ϧ��g-���;�ǵ����:���K�M:��:ruV����;��0��Jd���v�� |
�3<*�x!��v�bH
h����'ɛ^��
�1B����;�L	����|�-:/�h���W�]���M�z�`��q���9- ������Sᝳ����l	�i��zپ��3J8z�>ЦG�`P%8}	��%�޵���|�g֎�pR��k^A3�f:B�F1�9��˷uui�q:�k��.=�h%3	Һ�E]@�*��Qz��V)�:}.��$���J<n��7��2f#\��-�2�l�/0�J����|bcI��l��w�hm[!�!A}3&�tV��h�絯0%\�����@��Yٔ�긡,v�X��YE�	ΧR�yb���������(��|�G�m����3l	 A��cp���`�?'�OUr]uo%
� �攰�`lON��n��E?t1�"��͋�J �!���n�s�Q���꠹��ɑY�4�D1��x_�V*l	��3�!�#l����0O(%8��?�o[��>g���"� �bja����Ita�3��]Z���gy�b��nDmQ�>��(��p(��Yf��4�be��R�&��;P���������?(���O��&,��<�{yhN+����{�T���:,��}d:�C�~-�9ٕ1+3��(���'��.�M=��M��ӫ�����L:�\�4؏Ȫ0�9�D���I�H��A۾���`��+w1�>���f_��w��Y�葐�2����#�X�A�>�IN�8Ӱ��Z. 7dBbƃ����� ��/��8����X�s�R�|uu̕{-3�!EIfN<��^���T�Vpf����0���1}�e|lF��Xi��#^a��
��3��W�w�i`�(~GUd�6v�|��a$�4x��&���J�װ/�%u��i�0y�"�/%�M�ZT��=�ޢ�>��4�av�X�h̙����/��x��р�����3KE�Ξ�>�`1�Zj���}���3y�*YXP����g�� fj�,f���: >��{x�0w-�~���fl��Lג���]�7�M�1��N<��I�^��rOW
`�u��2_�ibk:r�^��{���HV���|�g��x5b)=i[�e��+��(�b�O�X��=�� �`r3�8�4�s�������P����uc�E�2�蠯���|� ͈P�ffI������:���M���(y���i�ڹŷ����;5f%(�H����|�}ū���[�����dj������*��M
dw��9��t�)�I��4��`;�p�;o�}�3�[���DDO�,�L�<�o2���6Bhr��-�o��s*~ �Y�g^�������A+�ƙ�Cx���P*KS邃=t0�y!/e���`��u����]6B���y��ǔ¹���2���JhY$���:���&}��F���ECy���1���k%W���v��}<�n{��Њ��ܳ��r8O���1Kͭ����f^��E�޺}�_��u�|��,�d9h۟ �AF�@�n�jf�Ё�<�}ʞ?�$#��*�%��Xyi��GF�&k8{��DL?��lve��J�JB�8k0�E�"!��I�o]����0I7[�J�5�1�fx�'�6I^S�ȣ�"��heS$Q����;EyQ,h�)>��RH �?Ĳ�slq>�1\Z+iЧǧ�Θ/����lK���R'��k�骯��>���R���i�C���$���k��{L��}]�p�̨~���I���$�У#�`��4;���}�Ƭ��+�Ϧg�\K)� �n�?|F6H��skobx�����krO�N�}*�bp�V���#��|�����h5�����*�-y0�(w܈7�z��m�J�>�/��͟�p�>G��[}}Ϋ�w�6�x?�w5Sӱ�_�8���X�|<�۰���t�T	��% �"KQ����QM���gB�Ǌ����$il}�Q��;��Y3XTE�(H"��y��;����ln'mH}h��[�H4��%������h\g&X?H1��s�N�?��VK��1�R��M����,e���~KjMsl�����c�{� ��ד��w7M�8���=�%�?��O����Yu�=��h&�(��í�P��|�N*�_#��F�/���*[�Q����r��}�I���nR�dG�[�d��QR�-|��_�
���%wT?���Zg��i���H��r8�o�ŗE���$Z�
)|m~C�b�FM�a	ey��&�-�t3Ƽ�ͻ Sm�@��^���i1̽i���1
�����e9��$vx-���B�ҥ�� �º�'0��3��]��k"U^V���r�/�����3V�6t�QHDb�v�o�HWc	����*tv���- l��t$����y�����1��"�����p����p�:�wy(�_��\�(�>�c��W�
��>z�G�Sa����y��d��S\=���P<ԜB�� �W�@0��@1����������
z4\k/��}kn�B�1&���n���2�L|���U �~:yW��>6�
yX�g�����!X���V�� ӻҙ��(�x���01^{���4�n�s���8=i�����ٛD=�v�zCH�*7���#D���YSj��袤�ɖK�F��hڛY�4��s�e��[����t�`��{ E������f��5a��Ibj�]s�O�p��\����sB%v�xu%�٦��ac@��+l����8,\?$��R���d����L���<�I�7���Ly��o̓P<�u�"�O6J����Q���~+�.���e���d?��mv7鮸��P�EZ�����"q���p�fS�)C%�Z�9s���"��*����#�U]Q�毙�[�r2���X\��̖g�٠����E.]��Կ	�nv2�T�}�Q�u�<�
����iɨ���I�C�Q�w����*§�a���P��Ľ'��|d�X��Wǝe�ډ���b��L2�� ��C�.
*bj�aB��-�T�1`U�n����=7�=�L���kS�0�L���VT���Bp�ӽ-����>��J*�݈�F�4JO�H�?����:	r`����Zh=U���<����{�&��y�O	�q-�Ύf�uݗ��/3�݇�:jb��EX�XU�H:R߽z��\�^#�z��7�=,S���"]�	¹�q�d���cJG'@�i�틌a�v�M�3�u���=��5��	����B�p��c��ŨK)��\a�.��4St�!~k�7�� I6F�RnҁEt'��/��{�]��v�Mm$o~��r��	��M�x�o	V /��MN���HW��Lg��k����J偼��
�J8�%��M��|kS�Ƽ&!�V�#1.��>	VvXbu��;���UcqՀ��a��/Z�A~��@g/+���m�R>��>۷��D׿]��7�7��H���<T��Lz���bs�H�J�&@O��tA�} ��d@8%��AJ��f�MNT�(@A>="m�v[N̼�&��k݀mf��^Y[�wsWa/�2�P�럧�Z[H�aoccY�r��P�_M�����a�� z�0�h.�=
e��˫�|~8�����f�`��ʴ��j��2+>ߚa$yVC����S�}i(��[k*=0יX��1z����F}z�p���7����愭Z�nw� *"NuR/�!�p�r���:��7M�����+��z���8�S
?�d]��ѱ�1���r��a�P���J�H�>������b7%A�J���o�wl�	V �����0	nX�$���z� ����3�����
�k<B<�UquO
y�'^"�[`;��C[0!믷Ya��w�K�P�C�	2�^��Js,�E�~f�"�+���x�;J�\�j)���S��]��"P�5�[s���H�Y�>�/��!�Qr\��-�J�u/����%�~�����
�3���|����޲lN��[�`��j���]ڍY�N�vϹ���:����em"�.�'�H�T�߹���?��o頌2n3�v�x�C�NU�R�]��l�E��8���.P٪�$���`_��'��f�!uĒ���Zy
�TW�f��V�mr�v���n�4����G�݆�������"��J�+�Ӽ�5�*�Y������hO��b�������Q����\���<��&��LzX�5�M����$����]e�t�����l��K���&�g�t�=6{6�5|����jiNd�Ў^A2�x������It,g�������o\Tko�:��lm*�U~�[ׂ��Ǒ��;��Q�6��S�2�r��5'���W�@��x�~���m�8'�(.�߀~/���&�M�3w����A���� )�`�t���ٖ�:
!�-�Ԉ����>�Ӭ�r[��. �"��Ͼ�{@P�ߩ���0�L��G����7�(V�y�%���v�!���c`E��b��@C�q��=X�Z�KY�W��&6;�D�V�T�*���q1�?/�в+)��;y{s&�~e�����mhv�B��H��)&�I#D!lP��>�Y�^2��sH���������W�{�A0r��j�}�Ҙ���.�2�!T���~�I�J�X�n=M5N��0�z+T1��Fmi&����������|Z=Lg��o~]�	�c���HE\����V�����U-�3��Y1��>b_���a�15���o��$����WI.�P�{h�L��3��C�����fRnR�K�(���dw;��OkH>���5��4���+�A{-`�|h��S�Ч�Kq�T��yo��|L.�T��3sκZX�8'� d�Wy�_g��*�j���}~��L3)ACh���\��������gM*�yز�
Ⱦ\m�o���#�C��-�ӝ�GqO��}�#ۋo�}�(�����SN���%P��7��W�����Q�zH�n���X�������>�3Y]{�1�h�4�3���x���Bƪ�%RF��;nM��a����c�,�Z�g5����R�sʞ��5�|�AmՂ(�&�%7��D��iկ�XHw�*��'��5�O��g�š}q��h�i�s��=�d�r�d���x �y��82@�OO�k�w�%��,b{��T:��R�"�ә��k�%=�l9`琖�v����";P�K����� 9,����L�0��&�q���a/#�L�!����ݫ�i�r�O	L"��T*��ޘ��O��<���y҆
k�� c��{),+DȬ@�x��:kϊ�����?pS����c枙\p&�'"����gS�-|Vn��<�NKT�uC3I=q�$����Bj�Z�A�̆N�+QaS6k��2&�YS��V#H����}��7I7"�������.�L�[ȿ�$��w���e��Q���`Ws�߅5"Ӝ3�F�!~��m`LH���Xl�B����_���~����ή{HqP޳�*�-: j�\Y�k.�1	�D�T�Ŧf���s�U(�'G�u>Q�I�-7�#�?V��u
HZ,��ܡ9�=a��AU���s�W�ʻ��U	\q�W�}�$, ��'O�M�7�U"A�V�H�?9ad�T��ź��9�T
Q��躄ͤtJ�V�i��cd�z���b �$z	d����v(N0�5OЄY�Q�K���Z`OJS�0�:i�N��̛�����?������Y1�q�rzȚ�1�0��v�#
^��	'��X�K����������Ojw�-B�T���AZ��o�_�AP�6xS�&�f�3��7�~�n�q!����g��Dh�p�}�,e���jh���;��X5����{��:��K�|�c;�g�z��ٷ�p��[w<f��Tt�"�놆��d��9k+ϱ
D�u��6	V\��QX��\�(i~>�VH��~���C:pvjR�=Ο,s�'E׮L���j�#�7�*�`���3W��Keh^l98��}�P�������l�2�_���,��N�{4��%T��|ܡÎ���N~5�)DN�9���@��R��&sCb��t��6Ǐ}����b\&R*��Ë����AH��fT�I@J��|��V��L�SI��q�ԉ'Ą.�kAx���8�*�dO5@�+l&D`�a����|µlN�YA%��u�W���xA�mK�mS���O��7bY�~)%ք�՘C%�q|O������%��2��(����^Z{o�'6��y��i}�����ې��ul;6@�k�.�T�.6o�nî���ҨY�t���5��9��n5[�Pƅ�)�q�y��"�Z��~��h�`
0�P�%�X���q��	n�쾈ځ�!�0z�D-����9�)�]Elwn�쪺b�6������ ǣi�:�cG�1�E�5.��ѱQ��_3���}�abj�p���$�t�'F�z���IH�,x�O�?��Z�}AZ�\���>o����U.���oyu?��zr�U�G�������E���p�!��W�ګhv&��J�h�s��H�ՅC��V��&��e�T�W|<(iO�Rtȩ1@�zŉ�~*�,��-{�tm��:����lu˻��|9�H�K�쉥����Aa�A� �g�D����zɁ���1�6�<�J�7g��L��;�	b(�(;�V���:/����������D�y��Ջ柖�{F>�O��b�&��7ū��v���]�7mj�%��	h���M�d�6�����T�DyG�#qc�B,F4R^|!.^5��۰�t;X��W#y2Н~�h�4ns<gK|�.a�·��ѯ8"L`&^|�w��K�.���y
P�=�����ÎF�3��w���49�p֖�Go����+�ܸ�E}\�Ks�u�=��MM{� v��-�+��n�
�j�-���	�b���pR�W֕�����}ЅeH�p,�偲?l�2��5����=^��yxL��U��_���x���;XYRo���~�]o`��$r���E�6B�L�~�;ĒWt4�#,s��Ӄ��p���=E?+u߽�?r�ݠ�Vu ��~Sp��y�9����fjX����B�3�`U~Fb�NO���@���H�{����9bS���{&�[�n���h�r�g
�<������T)[R��G��+'f��e✵ue���l�&9(8��J���)��>���m7�q��C�g3#[x0�����##��Tj ,�̠^��ו|Z�;"?d���Y\>n)ك�F�*z���R���*�{;��L�7�1l���iZY m�^[w�9$T��95���Af=�]�J̻G��i����﷔���XlxV64EB    fa00     8e0Ό6�"�M"ju�6Pg��>zL!a��b�$N'����?$V�{ ����DG�]����$�}���F�#"hQ��S��*}�jX�����`.a��E	��[����
�Rf�4��-�6�ǀs�࠷s���q#rN(����k��x]��i̻�3�Px���By�J�WJ>k�o���[9!έ8�F�!:��|�p���VY�Yz7�H�Q=,����4ѯ�CH�ԗk9�\V;j�� y�"kNu7������z�V�@�L2:y�{�x���D��0���Ch�HQ�^�z�0��J�]�1����f��g��<�&�ȕ�\+��(���!��Ȏ���MV���0��擭@]�[����CA�Kx �:a��g�.r'Lυ��+����LYcG	]Y�Z�^>��N�wu��mLF�v���cٻ_Wm�~��y��1���c�MĽ���}�|l�)+�&~�T'6��w�aK�<e�$�S6s�H�5~%`y������L�̆1��M��
�n����U�s�7�����vu��%�5I�r�xۼ��a���D��ɲK�KV��bƚy]{�˝'�Ahu+&*2.}"-���tm��4L�E� �xX?����$!�Jb��W����g�-�L���|��F p9�a�:�~�j�hj���H�o�p9�IX�	d�Mk��v��1�}i�6�U�XR�.����x��B��t7 �ksM!;^�fu2E�}n�z�'���V��6�yG��>2�O~��	zAr�#�ɂ�vuI���MŶ���؟2��98�h�L�Ͷ�2bU�2��/c�1JM譟�';�V�����;$B)W����AN����h��J��M� H����)q+P��:�K&*���gC�0��4qi�'��#�<�V&��ַ�x��E�aV��҈��^�;��XK���ё�K7lJ����'k�ڣ#�
B�18����~m�s;\d�{�?�ֻ��W �?hP��`��Dk%vC�Y7�����D���(��48ߵpy��R  �t*��,��.��I��%�s��y2�"�ۤpg7�2��"��XC�&A&d<ʇ���L�E�b�bmL��%�DE�J���T�u�Nj�/�(*�瑎��e:���h�X�U2V��#��f4o�����;���w4"��)������NB�Q�8_x���`����s�#,�4+o�'���r	�[{�CJ���2�����E�S�v�#b���g��)��_UÚ�I2�j ɑv[�� �,!����R�B�;b�g|i1����2�8�sd�c�9������% a����E�q Z���X���l9n���Q�[9���K6�Mz61�w�P3�lnc&�ާ�:h����k�DO�?�G�B��N�u8 �p��0H>ZJ���|ĉ���w���]�f��Ɵ��}z�9��������,`���x��Y�G�4�	�	J�SRkYbO�Vr&3b��[	y��,j>�/���Ʒ�5Ox&J��_�H&��0A��i1�Iܯ^g��,����Z���K��4u@���UJ������ 
�[�z�K�[y)��ӛˎfp- ����=�c̥\�I��]D`5��#O��at�9��MW�s���hXE�<��J�oyp�TR�X�"P,Y��攍�3�!�'�_��i6������g4��k� ��E�]���H�������6B�}ÑK�5]$����=]��=d0��+4��%<6B���"Q����@r>8;j���Z��,B���� �Ul|4�B����\�iٴڦb���r< ?(Y�=��n��ɡ�6���dr�]���n��+�Tt�CI���J���lR�~����3��Lq��i�؊�TK5Zg�f��xF�)��a}�{�`�a��� `���|$��l^p�L��I�I��ٌ�3O���U�8/���D��@N�a�rLQ�_;�����=ꁝ�_�͋��Q���K��~QiM]�������J�>.?Tw֪��DF3G�ҏ$,k�z�T3!ʹ��3ײ�"��'T�/���"��4IVقH��X��vێ�w��@��u�6�`wv8Qރ�8JG����+��o�� ���Ry�ڰ�C��V/Pz<v&E�x�u|=���<!i�-"yء�SŞ�Q#N]��]: z���ގւ!�}�H��tƄV㑬����8rqoFWd<`K�$U]��n�}*�/@�Oۥ��C'+#���$�!��JI�ɷP�XlxV64EB    fa00    1110Qљ
�&ԋ�Z0y�.�V!As�.;y��4���0O��ۯ��S)����+��Ъ�P�4��X(��y�9L�p���)����6�_��:�D��s$�7G�.J./�ы-J£7�n����ˤ�$]�v�
-���e��텫k=��O�)���.���w{{Ygs&&Q�p�y��ž���ݘ���	�g���%c�l��:m���4ؐ��*����r)�����C�,?����9(eȥn(Zm6�R����!5f��e�sP�̈́i��ȁ�g����M<�`.��R�����U���MT�>z}�:^uaD�P���\�D|C��!�x4b�P=#� A�y�����&��>;�GՎWi;�Y��fHL9���{Ҥ7��IO����V����&�����V]L��4�7�]E�o��V#��|lA����70�0,�}�q��L�[l���06�}�2~���3q��*��S��p8H��9l:�dqs�ݵF��pE�>A�7��^
�ʦ�F�u���׊@=����"]#�����LC���n��)p]Fh4*E�4@Tw��@1���oi����O)����t�j�Ƶ�=�1NsknKy��Z��3p��T(i1�������	�J���MSyF�y�E#�i��!�i ���`|#�V=��g|�Ղ�B��un^F�c��R�6|������\���⇹-y0$5�TC=�|�T$F�|-&�$�B�Dq�	6�C���"]�\�>�b1��}�ʇ��7�b�(�W�;ov,���ʛ~��n��0���6 �B\�4�)
���T��\W��/�FO2����R��#Iܡu&w��H������&H5�{�eբ����hv�ۿ]*�K�'a�͑�æ6+�$��3$��?J7��D])@ѥ��9��Hﬡ����?�l�n%����Wh��S� _�Ӻ�4c�|;:����;���֏�R��s����N�K ��}��5K�L���2괫��~����4q����ǹ��������������:���	QS�ǽ$����o�)m����1X�S���gɒq9�p��U)�Q�F��n�5;�8:���t�����c����)��88v��텮�nՆ/�N'#��+�哮��#�|ZFuf�sR��Vܶf��O��9��o��yI�F��20P�D·�x��~$�I� ��h.�r�]K��|D�澙��C
l����u:��{�Ix��sv�C�f2V�iO����uй���t���ᰐ^��W��kw۪�$6S!yLr�Í�a�
F>�K〱O+�"�4�'���O@,��O���{"/�,�/!6=�Ui�P�^j�~�W��4GК�o Q,N����Z>��s���%��X�ê'��Dd����e��A)�}߀�+��	��[� _�o�|��r�Zo��� �'�s���
�]�O �c�]^}��[]��e�٫��,L�ͳ�EDå>i��C��s��n��>ll��MtO$��~���8�R-�U<0�t�z%�MiyH�P���,]�~�n��'�Tn��b���!k���V9��^�h�O7S�DL���� ���iĊDc���~�i>
�\����7��QY��#��R.k �5�*Ֆ�sh�A#�dB�H9c�����p@	�UP� �_�5bD��������Gv��T�u�sŘ��������kj��Qd��ڶ�-�gF	:d�._�[���huS�gf�8�<5f�(
�����u�T��@��D8g�K�sh�MC�c�؍$�������X>1��T
}�6�Q�}��e8�'�� ��Cx���FU^��͖!gB!M�e�]�l����H鉉���]���^H���넶��G]z91��n �)�ցb�b��e�ܝb%%?��Sk���s�t��qM�,7�ŭr
_Ϊ�((\�����E��"� �t��ߟ��TIhO�ݟ�&Ħ--�4Sxf�{ Y"�w�������#"#n��f[�a���G/P}GY��q��+���w��0e|�.�^ʹz�HCg���t�)�ԓ�fG�:|�⾅��x1r-x-%(e�~����I�l�T���8������
.e>���,Ύ/�~�ʿB2ه����N1s�`�9���"7t2� Nh�1��:���=Ķ�l�u�q�."8-�)k2fb�g�sj }�M�#�Q������7���c��<��؋��4�Eĝ �����&Ю��\&TC�m�Y��<�f7�R�:�U(QK���X��At{��ؙ��1��bq�I�'OoA�B��ඌ�˧'�U��r��o^�����jS�+m�P�A���x�m�nK�<
������[�@��g�Y
��b�ģ)��;�}%zy+�Z�K����9QU�S�KЊQ.���}���ax�b�4R�w{�Y�$��i�	t�Nۇ
X�cѣ$w?r�p�2&IwW�G�I�޷q�����sĢAL_W6@�Ɵ����v�8�Iv�-�@
�9^��F��5�����O*�>O�9�W��T��D��"@6c'^�LPJa�{���y=�+��4)��k�z����xĀ�o	3��!A�o���&׬�
J�|k�4Z��R��Q\=i�͕��}YV����HY
W�-`���7v����"�6<�zT6d>M��^�"�T�@���I�N�x
p;>���m�BBV=�����|�N3��@����~�I��.��*��%�腿^$��n�ܯ>n�;)�o8��c�ډS#m�ā���붩�$�u��x��$C�u�G�s��@z�/d�
t�%�o6���F�ɝ������دc�aqڈsF]��L&3`cj�7�د>����:5��,���oҘc%�`��/Xb��4C�3��"�T���?��-����\���O�NpK�@��43�?���n�W��er�j�V�,3�|�Z��S{��
U����f'�[T�8f�Q�:�n�D�~\?���4,E��)SSHݦ~��[��g���N�����~�ԝTa�FJ�/˛G �����T����杺cO�x4��H&U��K�$�yW05��wu�|���Fo�N.���W@��`�Z1t#�:�8����������(��r�Èi�A��P�Q�V�YmK��������2x��m�D��ݙ��2�*}�\!ZM�FK8(^���:��~97kj��.X)�����
�����io�ϟ{hz2h����ʨH�0v�.J~ ��;Ζզ�S}QgΖ�o��3R:ڮ1C3�8���6��R&�P��>_�B��u�P&�\���l9Y|�;}T�u�N�A�� �-��N��$+�ҜWw���t�a�3�Jx_
QRz�At�Ω`>nxV~:��vt��pLX��T�b[z��R�6�}�]f�G�b3������4ĻKeY]�R
c�����F�q�)�D>�]/�y~1��7:��׮3z�\�#��r*L_�)>A��֘�G|�3���� w
I�(��=M��"����Vcr�3*g6�g0��p�x>ؠ#���B���-�B!a3��f)�D���1�LG0�Qm|
ٕ�/�KUő'�rJi���(���DO7v��h�K�lb�c��\��� c?�.F\�+B�Eޏ�l����y��א-ĥ���;cpJ!���z��C��!r+o���yC!�L^;��	��i������{��������ғ� �V�Ip�L�+$�C�hV��ʂ����X��G��	�}.��n�9o��W��ӽ0EPQ`+�n�1�Z�V� ��{F���[�6������4�0���V�� ����\��[����b0��w+͊�Q�ri�ғi�|�s�C"�������4'��3���a�8\=����PG���&��ɹ|ɸ����tj��"���^0%� 0�0�>�*���@_��7m*��SU�QK��sxCUND����`$�ty�����NET�F��i�⿼�&�=��i��h�f�5�9M��4����Cqn{�$CY��S6mc��?&0[��~��n ��^��E&v)�h��E�۩���]�����xAU�%��@'L�yT��/�X���&��fH
�SN�JO`�A��ה����s�:߷t$��/��d[0��o�Y�k�����kQ�����WFp�N��]�3cqx�z�ݟ��U�)|�1���?*��HN�G�w���i��u�@����B7�A�OH�O�-6���~6��kp�g�? ��m�U��.&M�Q�Vf�Ri��sV�"�X0�����6��H�wXlxV64EB    fa00     ca0$-;\񧟾-�oP�BQ���-�;��$%�aj'�au_��v����^E���x8'��X:yĊ�v�+�C:Ƽ�cƅ)%���t���w�	t�?���p�m��f�q�2�VZ�w���n����c?4�1���䔰�N*-&HS5Bg�HQC�GSYnJ��M���kͽZ�*�U\�>�4� ���)k� �E��T��aĢ1�aL��e���n��$K:�ɉߩ1��g`�Q5�L4za����x�/A���@|b�3��Ô���^;�i����&�9�WWl�S����N�&�:C�%���p�	6۫�s�~�5/O�R)˨�}��Ht,�������j����)�L�~��+�/��m�H����)���/�{��1�f�L�V��5Ȍ$�eS�R���r�w�y_��\�%^�E4��iA���Y��wHg���D"8p�c�!�e���Xdt�z$��2ᾧ�>��i�N�f�q�Ƽf5��Jm���v�`l^(��E�4��Lۈ�iLlJ(Nǌ�jO��^ӾX��"Yҵdj�(R�&*�ڛT �ga�߰���YL]�^�y�L�K�b��";�9K�%��'��������$����j�c��Ƴ<�v��d����ϰ.ba0y?[���:����Zp��KY���RG��y�<��t���WHY�e���媏	���X�\��:ȑ�Z1��(B���**��%@(�ί��������m��ک��0���G���f��a"� ����D�������/M��"|��"�U�r�7��� �J8����%&	��]>S[�B�;��)`�)��t��x��A�>�ڴo��ޱd�*]nG�Hc��nP��(�2v���;꺔rn�^cĘ�I�r:�X��)�����c�jxt̻� �R��?��jÊ O��I��o� ��.�l��ٛ-Ӏ�qL:��8yA�3���?�nj ����J��k��hr���n��]T�U�HR���-/=j@|[���>�^L����a�"i����1�9�N$W�,(����vx�e�*G��z���#�l��}��To�b�������u��<�o��AK���<���;v���m���<�?�`e!�x�{���3��-�&b�G�x����Q���^�t����,yoҶ(�<���Q?������(�6Lszn����*��Dk-r�Z�K]��I7���'t$@���m8�
9IL�g%���R�c P����e+��:jS��6��YO�.Q���^�<��2a�N��f���Y[�֛�yI���u�:��6t��eys[)������_m,����Xx�X�ف���C
2(n�FJqچ{)~�I?F#�3n�m�m���3�߆ d�{G�i��
��#���7��>����9�� ���Xq�ԏ�B�+_�3C,"xS#jl*@�3�e�4���S7x�9xT#���{ɣv�F������@S��5]��d�����m6�T:��i�ѨX����#n�n�У&	�o����T���!���l���]ʔS��#�G�rs`��F��y9ɹ��L �
�j�t�P�����ٱ�?�"�W+:�vfL��}Ӫ�cf �ģ����C`9�7fV��gɰT���!��[����"�r*n��|k쑧n� "a^�Z��:�"3�F���I/�s���6.w��֔P���
8���N���R�_�%Iش��|���ZO�\�y�GuaX�Rϣrrp�/+�B�Ypw�������D�^���I��瑘X�VKlh����S��	�b����L�{y��Q�(�h''�I�m&�&UiԀ���~��y�͞�p��`�ߞ��T��M>��"6d%Y�w�q�M�)DLZ#�H�cÝmk�v��7ly�>PN5�G�O[�J�������-��oa��Q
Ǽ��fSf�9��+$��҈�����y���v����NLd��S3�[<��B����R�J�8�T��S�*Gp�Nd�3|��s�{��\`j�_RV%8-�m?�6P�^^����f�`��P{g��+��L��L��}6:�C����'[���^e�ӡ>��3[�hMx�+@�6�YMi�az��q(�{��avbF��#t_�6�����-��:�08���}|y�#lz�:�w	cj`C���a��q���b��qۘ��1�A�ޔ\�z7�f��'�}H�?���n�O�7��XO\�E�tԺ�޶B�%�o��jJ��׆i������ꔐ�@Y{��	�)R`�gN�ZNp���ά`~�?�ي��D3͋�6[������V��v�<M9Cc�<����o
��ֺ���<��[U�r#6�y!FF�=���i�>��6��Ua�#���4W�FS4��;D&^����]	��A#p�J��1�x�7%�0K7�[�=��.8
3��{�6p���՚�^��!�d�tb�B �TW� ]�km��ǭ����-��c�jU��T�8w��y��i}3U�j��m�T�~�p�|C�&�����D�E�Fn�����^�[�lV  B��M	�W�Pp&�Mj��n����`j�
�����D�&�w���lae*dM^�Q�;��E���˥�
�#+=�Y���%�� ��3O�T�`�<��3�P����ù"Y���)6��2�H
����R%�y�5��q�_����1�}����=�}��ok��Z�֍���Z�mY��'Z�lC}Lz��Vh	���bc�g&��po��C��Bm����W�*��X�����[� ��Q��l��Ρ�ۊU��AD,n���������'Cԇ6����*~
�z�vY{�u�UB!���y�i�7�)�"!?������(0��3�f�f�w�����N�Hw��!�L��=����b�B\;dP ���e���r�t�x,�f.8'����=3�;9�w�B�ۇ[����i���d����aq#��i�ZeC����e:�)�}�OA����	��d��!�� a�}�v���T2u:�a̢7��b3�FD�.r��Ѹ��vc��[[PU�q}A{�:Wbn��KQ�TT�z��>��ܤ!~S~�:&�+�� �
�zBKÊ�?jeQ�CE^���L̮3V���i:p'��O �\9�2떧	�-��x���=$���$����[�����/�J��|�i���Q�*�o�'P�N����L��XlxV64EB    fa00     3f0]n�bLEL���������0&������ ���2��䱐�f�%)u��q߬�7"�Xrך��i8ÿ��r�u)���ܿ�.q�抚}�[C̼�8X�6�D��&6�#�A]r��F9ŕ9���9�E�;8NP�|+^�A2����P���;���`?r&���"��F���@�O�N�H)�v��P���)]�ȇ����<� �.����l0�xu	�:�1k�0�4��u�~`)��|�lUS�o����VQ�B�d�$�xw�u�!���s�Ӯ���d��:���ڒ��:uY�'��W
����i��#e��EU�Uz ��"�x�Rn��cK�va�h�$Y�_�}ne���H�B��6�ϕ�N�2cI�-����~�	b?�|�v$��̋�Z�A�zc��n�]#Lu��!Rb��9��!��?���c��3�;���p,����&�DF+�[a��ĸ�ȁ��\�fy��G�7�o&I=�7)������YF�L��[�R=���UA(�T��cF�񰁨.�	SgГ�wa�
�3l���v]�߅���{�x_.�Ѵ[Wb��	9�bn�!��!�0E��u�.FH�~Ã*�һ�@o{��e�[R�����6��@�lः��oԋx<�-(��;Jk��!��6Ey>��U��Y+ ?/B�ɘ1���l$Ȇ�.y�]$�>Eq�;pi|�a}6����3|�t�@!�D��
uJ��7� ��~��X�q�B25V���d�T�׀�5��߸���:?�eq"��j��r�O*��pgY��
��;�T������/�^肀$�ކ�?��"O����>�K�� �?�F�m13.���qM�84t'�̣�p��x^�����s��F,T�O]aT���	'?�����͎EX����۩RK��71���n��\�մ[��r�e�7�x�׉KQ3�����M��2\MO�	qsu�Y�+�K�:R��M��=��rBy��L��XlxV64EB    8095     b20�K,�Om�]��<ͩ�⌓�k L�	�}Xc�&n��<ӰAG�w+(��K4��@���0�*��vc⟈t���Ȭ�5҄���a��ݘ���K�&Q�\��{���~ h��.���H��G�F���2ᱠ'Z��>�:�Z��ʶ�o۫�=5�p��6�l��Ę�Дd\ש��\هXR�g^�{��k��(l�l�4M�^+7ָ�kJ@K���xU���\x�"Op�͵�|i��dU��t7���	����-g-���C�����]������5��#���{��3e����^!{�j߄�Av+�u-��E�6�F���}��C��R`�?�1���q琜���x&X L�!��x�㭖:�K�hjqB�'L�TW�J��KbX.�����'8�z�Q�"^��h_���? 8*۾e� ���� r��dNp������vJܹP�8�Ԯ�>���3�(�ob�X-�gr�4˴��X����봗ʤ�R�F.���a�NV8x%���:[|1�K[�Fe���g��.���B&�Y~�����p����נkS"��]�f��h�����Jof�~t,BY�6�;�3{TI�FG^��N'
�TA�G�4���U{��n��p1��N79�+D��M��T\ ~s8g�2P���ٻ��w��&��</�n��b|�|�A��
6B��f��Y�)�\}G���hMҽ�ؤН�-�JV��Q�xp���gfk�#s_~��FR�����������~�*,���&���8ldQ��6�#)*>R���92�4�r2#���N
VS����^3����{��܇�$��~�3	רּ�Xx=vPc���F�a�,��:�Ʒ�h�A�i_�i�s!2c�Q�=싊���O�����tj��Z#f�]�O�,wx7z�*ʾ��9��)s��ST���_����z�����.\ɉ���=��,��^�H�#�7��Hy�"B�eM�,'���ʢ����&�ǳ/_j3�`�rp����}9�_.���=f�@�ʂ��Ft�n���]Z�64��S�r�J/2�K�*���4q���]���y����s�wH��9�8�0�SR�5����|8$�Q��/�eb�B��#g�-��m�L����ֲ_~������k����Q9᪗Ό3�/p ��s1�?�K6}("���Z��cn"��5@&�uAΟ��W����j~h(���5|��V�R�P�+���uAf��R�}��PS0�[Tq7eaa:��C���"3��crn�%r��w�o ��tF;e��V���/e~避�V���c	�={7v.{��;[P�E�x9P0��q��㟢�z��^�yм�UAɻJi�vY����	d|�M���J�Cz �8 �Џ�3V]B��!{�ǐ�Ϟܩ��*f7����d�8 3�cI$���op��}���cwi��;�*��p���m�V��9�u{��<l�j�9�N8A�q�֛~�V�_!�|�e�f�W�@>��Q3��
����l{_����!*;/�@4�����N�z��#��.S��[��|߬����H��#��ĘI��a��@_K�@M-�EUOW�Z����]�3qwGX��
,7O5����;�
ː}2a����0yɅb56���l���2���_U��b��2O��
���8<v55�}a�d�f��m @�ű�ir��W���m:d;<���!=ZD��	�x�I�PɛfU���[����:���S�|��;��;$�2�NҊ:?n]���q3��|�+�Nb�lb�擰1ճ:�� �$&�y�Ӌ'F���F�$B��%�[X���E;��b2��@g���F77?X���[�o7o��e1u�;0��Lx���F�) ����׭��)��~w1�!]��L��"�O�Y��%*_��ٙ��f�*pg<Erl쫪DW�G�Հu1^U4B�_��I�<��1qT������*�)���è����Sj�x��Gw���t!�.!��o���Q���K¨��GQ�f�-��hG�)2�j�ꛓ�K��*�~�̙����ё��>���O�,�P��)T�&^>�I��V���d�v��k�:��"+{�{���ܕ���7�D������x��]��M��0��XxQ�Pl!�^뫰�Gs�B�c '��LL�.������.v�C�gX�>�O_���H7ģ�;����y�N�D��o.�c>�r5�C���o�k��T��Q��v��9'��X�+�6Ȅ�����~��U����n&8�/б5��D�0�b��-`MY��`Y7�6��;�M��6�C���9����*y#+��;�9���Fn���ގ���[�ӳ�R5v3�Y���O�}��Hݳ�j��c?����W��s�x�)�8X�'FǹOO���s��G�����l���AZG�:6Ԡ&�θ[�-�.~j���!���P�#���T߉�x7[i����,��^�qVʾ<S>��2A�;'}az���sߟ�
q(���w�ז-�X��9�TQ�u�p��e%^�F&α0!��:4e*��&��Z�5�\������J��Xԫ9�!����׸�O�x�������%�W
1�!|$� ,���=kS�u\�h�/�b�KMpG;�aѢ��PF8K�@ _��%�[o�iwC�(\��*��RN�v��BjZE8���eHgJ�ᡮ���crE|MD�U�����o��$6����g��KSZ&�8�v�;旃���);s�'&���^�xK� �G�p���h�a��S`Sghz3�&�����-=��r�b1��;7