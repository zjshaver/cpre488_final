XlxV64EB    5223    17400C�� ���
�5��%-��[c#��@	�i��#��dG��!����H]-e��W*>�X% �nn.��J�Z������9�� �t�T�.Bu��'i!\��$�K����/�&uT|ƿ2��#ǆ����Ė��Du$t��s��;c�*=3���`�����5o��+q��i��z,�zU| +~�uݚ�*6��92�b�]����}&!�`^Z���^�;������눜.uk��CH\��:R�[j`�������\2Tٚ���5�8���ӹS��Dq�Z=�	�T�Vz/B��3s6�x�����{����{���"`Ѻ�|0T�hD8{^���'�����E���D�F��~KN�a.�٨���u��J��Qm/�>Pp`M>�6_ΥP%�m85�MOE^����3<�^/�����4�/l�h�ΥL�.
k�O̕�r�b<>pO:M�ؾ��M�h-���w���n�`���$gH�j;�w8�#	���~R��I�`HI�Vo�S�� �Є�Iu�
���s]oj��`<�>Ȓ��Iۤ�F&�5�BSPE2D�g�� C��/H[��-�䟤[
�`
�k5�P2k�Uy�Q*kXp0b��?�[	V����G�.�#=k�co�e��K
Q�=ه�����d;�k�2#�����e
(�w��#�^�2�Y�;���oA�f��a�a��f��H�s�NT��*|c�#�� 2'�E���וညo�ϸ]���eSy��:�Vdw��]����p����#�g��
z�V��T��
��ި���=���I5&���AQCKÕ�eQ�s~1��g욊惛�g]�&�Jui�o�z��񣢣��%͙�`�y���m�og�,��P�;Ɨ\Z�#�9)-x��s
"9�WKZ_��%�C���0��)�$s��DLnǛ(��AR��Oh��	����SR�J����Z�f�� K须�?%�oAg��G#G��j��Z���?BuI���q�Q��CA�^wv�E`26���ԉ������͉��Am�l@����vDAmm\��J[`j{�  �{-�ov�/o���$�(G���P��4�V#&ܞU�l���
�c��Jj&��óņ���D�!%���3��}�.G��0�	�V4�A���q����n4�o�<�HD�ڥ<�a���Ήy�i!v?���l�	Q�����i|e�����p4 �	2쮱���رԴ�I�,�މ��o��i/�qM��\ �V-z$`b�l�JWf�f��
��ڵN}~�[�7����Ç�G�0�1m��g��KZ[��bg�W�Q���5��<���K�=eFV#5� �K�~(;
d�Y�P�y��#�\�f��ɽ�u���0+�p�ߥ����H�I3�ntw��fk�i��Yґt��	tt���6���;��+�eA��4̟�!L:��W��.�d~[�^�b�ef����X ��\|�̷�/��l@�T��mVXK��-q�����P���_�f�Z*���4��M�N���#d��%k����9����M��Y�)	��s��4;�nH3�W�:��=dd����r�$[�]I	�->?p�8|4��1�a*;B�Ya��A�r�A�A�ۋ�BZ#m4mgb2"��R��㖣��oa�}(ӯ��(T��X�A��8�c�]�hH���&8ބqw�p%s�u�(�&����\ ~j��\-��>&��&�7�M�㴩���$thTb���t���hY�-CŦG�X�{��Q�]��)�F��f�6��W�����X�t�Ĵ���Tt���V%v��rIY��-&��b-F#�P�A>��0��'K�H|i1���uŁ�HVԍ9a�Ƭ���E�ﰓ�ǧ���";�SN�we �[L�W�:Ɗ�@���MP����-�������/h��6�����w��d�gV���[S��Н�@�>��_����!���#�� �o��)����xp�����[?��pId��Mh��ͼ���H������H��WLFSǓ�1�#�~ӫ������'%p�)t`��R߰�W��"�X焤�� �r��w� O�.���4.�e�b�aTR�k���`� ڨb�N�
9�+���̘X�����{��7��R �3Ez���qԚ�wm�LxCD������t�ϐ$LU�dV1 ~�����T2�|�]���܅��L����+H>;���6Μ�9�5�Z�˫�e���]Ϣ����Ϭ�?.��&��޹.&Dɪ$c
��襥���W۝�:��N$ݹK�>
C�#{��pM���kK�)p�H��z�X���I3��n�cn�?�e� �_��?�l�4���vu���QN;�i�"`�6�t�a�l�����Z�#!t�Jt> {&�J.�8~8����+�(��8��>kJE��JJQtND�8 �u���A�����0_�A�d�Ȝoô�?����Ef�OfQ6������7k�M/���Zt3�N�lDZ� �͂��R{�C��c}��x/�kd�ZYXQ�u�~�@�c�f��,?9�\���7��9�+�wY��M��Fx}j��q
�9J����-�ܰ���~��7�2��8�3Z�g�Ӹ�I�'s���Zz���I
�4!ZF�_h�)��XDݹ�#�(u��^���� 9�AYL,3v��,x������1F?C8`%ΞR=�-�]�kB���D��y����>�'�UV@�z��,:��r��id=�l\"����.��`GJ� n��b�B3������Jq��S"��<���0���z|�,������*9+��3꺙�<��U��Q���=���U/�/P�N�!��>�kQ�i��\�&���p�إMD)�˦҇j��%ɋqΤ�5<���K��]v�>;_񃔃g]����I9��xƉ��N�݄� ���M���ph��Ī>���4�Y;�V�y��3�|��bO���#���#��a����_��%��c�1S��G���`�)8���mM�)��O�^0y�"�)F��{��&���D�y�{�O�>�.���?�I�M�c�_�{�[�U�$}|��"��q��P��x������2���2ymX�J��,�u��\@���s�yϐm�Jk�HN�2�l��2|Kk��|��,ƴ�*٪.)@b�-�A�E1A2:���W� �������(4Piy3!�X��Z� I}Xs����㻸� �=7�JKXt+�7��t�k}(,Zh���3`/�`��H�X~�6�}�k�\U�cH!�1��\�U���W��M�����©���y����ટ�Hu��K���0Y�&H6�&���2/���C,��g3���%ǿj�
�賁x`E1�^�x�<���s}!k����>�s�y'PHvͲg��H`Q�s̒���t=�����U5�+�l|�hA�A{My�|�⬚�����&bT㹮����J�3�ۭ��(;�K�>��|I�ϩ��[��sM�!Ʈ�l�2�z�"�����H���
�����8�mڵ���B ��r�C��y�Koq�ܥ��.��r�{Z�E\1���_y�}�zo�Iʥ`u�'/,�	�L3O-���B�����5w5�F��`ٺI�2�������zI&Qt 	}��&X�5|U��EM�����f�LF��F�����3���[μ3k���.�!������i�u'�fW�5|.�C���nBk1#`M�2��\����!dی!�)�l!�
��㊥�.$9y���[��ߤ`c�H��%8�tď�(��K|I�ǽ#��j^֝5t��f1�.�M'n�,���w�j������"0�/���B�D����A��bN��3)�'�ぽњ��6Qع$O�p��2理P���y%yo�%�v�)�?5	f��:r@�Z�2Rt���҆�a)�K��� ����x��&��8�����(K�"�$Y軁	�;�;[�5��@��P��r~��u��I��lnA�HB�>�*!��*��*F��89dZ�6"]�%4�r+[Qgd�ǋg�lѽz�LST��9�ԓ�*���~Η��֨�e�".��6>���b�������-q��<�ʫ�W��4�LTc*@�js�#/v�xw�OX��C��e��c
9���E������+��~HrR7�FP�����%�՝��PZ#|Þ]0G���G9>�O�;y>Z(�k&��׳	WW����xf�����+R �O�x>�;8�-�[pB�z���n�����"0QË�w!��*�4n,T�S��{4��6�v��l0֢����V�yВj�0�F���Ik^7kC�y�����̡�w������/9\Q�
�O:�1��ͅ��H�]���� �(�Cl^Ş&Z�;!.`Q�Ӄ�dh�W �^���h�����w���#Ŝ�dɋ�虿��`�>�A��k��-Ƃ5n�1��m�|�[O��̓n%��po+p�-d��u�-A�.[�s("v�e�	1�m�$΢��g�QZFG�Vr�ƭ[X���a��y�7�rE�sw��{h�?��z@1��^�G����|���o`��㩦���{�;��A����>�ጆFCD@�1���q&�%Vur��e��w�V[a�ap��$q�̳�'��X<(��{�\3�G �z����_//�y[�S���%��������2�(�~�_�+���V'��~���`�,��S�&qr\���:e�P�b��D/}ي� �ص~�g����'O�p@�*p3�ݢ	�b>�}5���f����Fa �?����v�����Ł��	��+�̖�S�N��H�����;��2���l����`�>�������7-�"j�K?w��3�h�9���܌.��cB�{�g;J+^4�:F�ʺ�j��?��	@��&rnZd��zG������<iɛ�A]0{��;Й�P�����g�G.O�6���S!o����9}?�3b�+Ǔr�D�I��1ϓn隐��[�3�[u�81D�)��& �����L�Ur��
�\e"n�7��c9�V�fQЇ�ԨLשV�	���X	�b����4Q?Q6R��(3fW<�:o��v�Q�#̜�CY���6ݫ��y/����d���(Lo�h��y�t�z�}HH�AeS��	i����a���.��.	�WA�D+o���bܛ3y�~�����l���Z]�a�1w.4�.�YJ�A}m�|ŵ-5Yȧ�
I49R���?�I��(���p3���v�
CMhFA����o&<�����H3\S�T�@���R�VKDs�%u�Y��5f�t�,�P?�r��fFr�j1��}�liM����Eb M Z8=~ɜP�r|u�(C�(Ne�A}�UB��ܥT��0kyZrH���g(��m��Dc��IĎ=�������Ϝ¼�M����rT_�;���JYNEw��)��}�ʚ��>�Cǂ��������ñ��l��b�"heg¶vVgU��\>���,����\y������or2��nѨ�؞�8-d&� g����� 	*�%�y�[���ˣ�n^W��/Uf�DvSQ���(��R�����o��I��#�*g
�6S 줳��b�rO/�|n�34�S!�[`h�YԲ�5�<Õ��]��"��HD
M>(����w����\zE8^'�����Z{ ��3��>�q�o)�Ta�Q㑨���8}�� ��y�
'W�OL̆�`�#>�_���S�k�"�1�g�iP�����������^��ЧE[a�N��D�.��WI�~pTO�!��-	(c�	�|L���AJ�&k��<j@�I�����erַPYv���B�������Ǒ�#���M��!K�vE�k������@�i|]X
�`�lE?[�:H�E�
~f-=�@�R���D�f�h?��