XlxV64EB    b086    2540��ठ��8���t�7����X�/#l�m!��?〴U!���1%�r���r�.��c�i�jGؙpt�F���٣*�b��9pd��:)��H-R�B�8�m���Bn�SK�_� �����Si�E�3��^�,�k��;�J�_��M@����71�1��p���b�N'�¨����zk��I�Œ�X`}�Q+kD@N�sո��?Ʊ|�d�-U���k�I��[q.G��z�����X�Kv�;�}���|I�D�]�:F ?���t9%��"8�4�?5�r_��xW�S#$��}�����U:�F@IM�r���Q=u��?��	��@:9T�h�%f��� �T�����\���i��n�ԑ�7�V1=>�8IfǂG�'�xDc݄�ب�H����P�
}�c�>ܕO�*��y�ƅuˆŹE������)h똻�2���*?�lKQv��c�6�^D���;��Y��hX��&<�X(xy�'��r��d���,����0���F  l;j�����q/�����W1۶:��Lz��p-�e��2�3�d@��cE��b�x*�복B�9��T��|���}�{��8�?�Ӳ_���٢~���I<�&��n?l��<X��]fB(=梦(��ja���[���ww����sV,���>��ߘYtAw�M5��܇ز��&Py��H܁�X�����
�s^�X���C��3�2�Sh�j�xE�P�N���k��������Nʇ���d�Q�.����9��V�ř� ]����d��qe]c'�P��:B�hQ��K
�,��df�?��ګv�,������T�1�%p����{^��! �Xw4}��h�A��a?���ȑM1�u2��]vU��!i }	a���beK��j�Y
�"�D����T�B��s�\ÞR���浖T�'�nY������O��'��y��HN�t����� &�4��=%3D�d�^�@@���I
����� Fߎ��pm���r��zlH�K�5�q�2;��I��k�c	0x�/��:�8��BqX����'~xC�F� ��K׊�����c-���[��_Xi (#�/���4�
���}w&�f Vk��KG���QN�>��E��<c�Tbz� 	�)x5M
d
��0�+R麍v�
>r�d�5X
��
��K��=Ġ撂9��j@	���hGOd����q�`�P��< ��!.��IWB�����*]N�gɕ�.cY��='�0=<��CA�*�xdh>�"{�Ȋ�t�c4�G"NQ�(��V�2P��*��\4�
�z�9^Ԗ�r�L�.B_���d���!Å��Z��@eH� �W����0���
q�Ęͦۺ�[$Y�}����=/�n1|���@��\�xʹLk}���݆F8��_ǁw��xR���~ߍ&���*C����m��µ4�)�'�[6�����p`�ddV7�$�k�դ*_{-��~Z� �/8>!DF�ع~���Q�U�Ș�B٭��ʁ\y��pҌ�?���:U"�fa���}rO_kuJo�ԍ��.-���9H-";�p���N9�'3�s��v��\O��,
J���1�~��5� C���'j�MC���`�{D��淃�ShR8�
0 n��D�<F<�g��`r"zj ~>����퀍_���c���O�z�,1 ���7�TvR��<bc'��E�n^�U�i�]o��?��1W�͞�A��j�M������#�F� 8���d�3�yF����G0d����@���s��=ף#���ױ+/�X�P:θއ����p�^>�,�g�K� ��:A�6-=�,�m��mz򢨏Z>�"�ȿ����n��iQ۽�B]�%�eF\.W3V�9��{b�j7�a.���8��9�q���!�_y{*����p��|����w�B��t!��,�2�@��&PF�B/;-#Z5���$v����4��`�'p��� ��O�ef���~�5�RGB�=����4#Z�e���4����(U}�5B���B�E[M�5��j �~<��-���Y�W &�o!}��ɘ5V��ߓ}�ר�����#/[X�7M?��c� $�jz�̊�x�.#�&�+Z&}�g7�>h�c�`�%��X�{{�/1Wcp���1��6�D�$�ٱ��~���ep��L'�r�P
��'J�_R�@y[���e�A�7�o94��d�����U��v�"N�&(�4j7�"]���.�[�@��7_^P��!��L�_�2i<���bM�"���  '��tC;�Ш��X��#}�ng+̡3��b1�s{Dk�p!7�i#u?~f
0��<�x]U�@�u�f�v��ͯ�wtT�c�4>#����S@��wgn<�EG���_H`͂ /%���͡��<3��՝&�N��h��WR�q =)���G�?M�S-�o"�o����>������{�7�?$T�.oM�Ⱦ���,h�(Oo��'�1h6��[���0x�������sm"/�X�g-���|djc�	�6�,�9���ZG�����d���X���1��U���n�k��RO(��7���H���y��p�F�{�'I��4���S&���[|C��oL[Z?Z�d�}�j��+���Q�^����/���hr�~�kOX}��Y���{4���G�B-��:��.ߍ�C�B���a�N���x�o�9����~Ew�q�Jڳ������F��aU��Q��b�o�`9�A!��B����´A�M�'�Ċ��t�B��y�x�k}�"�И���q���057��E�;*3�ZJ0r���I,�������Uy1���<f#}�H��h,C.2⑰Q��#Un��M��-�R@��������> ǫ�B��7��,�����j������*.�e�����4x <������5<^��B��Bnx3�V�t�g�O?8x���� �l>Лq�����.�������Aw�G��f�.|�r�7!_O:q�RG�Ǳ6����?�Xr��e@���&�@s�x�8ـ=��.��/�d��t�]1T�Su��@��f���_�:(���V"�f��p$ ��(g��肈H�1.��yOCi����_}������G2�Q�,\��8!C���򥗞o�$5
��;���f>f�Z�O����NE������,�2��~MGX�_fD`��7��jk?�ӡ�.r$k��J�hqeΝ��=�n�3�+G.���q������C&��)iI1*.�.l6�EN����_b���S0c������ll;]��N���4��{�;_t���I;:�g�Ú��{zփ��>�F&b��v$<D@Ʉd)57���΁��E	/*<����b� ��a���xf$��"-H��iP�o���B� ���8�R1*!��p�-�R�G~���(T:��$���:�s����A�4��^�TNF(��`���kAS���"R4=���Rc�aw=����y�G��i1p��D�n"��h����Q[H����'aI��"P_ya9	�Ĝ.}������5���'Ӊ&!|��&a�G��ß���I�_�C��)��Ȩ�=�I�#�^Ի]+-p���Ed�k�d�h@��g٫K?���jY�@#İ֢�`bp!���F��t~0&6YON.o�.��hh:�ӭa�c_Ee�ā8�5�ڻ$ml'ճ���&�-|D^�h�oI$�շ���Un�	�Y[����kD?�EΧz���+{N9/,}�^}��8��T�3}���oN}&�n�a,.��kn����3F���;�u�Z�'�Q�r�T	S����×�@�F��,�f�ʙ_���f���HE$�؝�{T��A�!����7Ekr�t��D?s��zosd��V�R��]��E���pV���@aJ���q��J��%���|<�]�~L�;\�N$���T�U�R�h,�1f �k��nb�BI��$bA/۠JanN� v� ��rr�!�A��m0�Ы%�*��i��^n�2�$�j6��H1`�C�����p���^������t
�����o�������D����tk�ƺ��`��Y�ș�`?��y�#��oDH���-cg�i�Jm9������c�#���}t�r̬��f �C��C�V�ɧ����n�E�N���v$�	�r\�-3ӫ����� ����	���X�xQZ�XԷ��`'�z��iT�>��[��ε�F��R��fٌ�SE͌^���"͌�=�WW�>%��y�|5\gBR��i�-�$�uS��A�b��5��I�HUa�(ܝ[�UE�|J�j�i�͊d1B�O�:0p���+I���z�	{
+TUN" b[.-�!Jo�W�㞫n���v�A�3��|2���  ����Vd猫�8%�0�����oʽ46it�f
�i��3��d�ug/�L�Kz,��J���M x��	5|����We�'��W�kkL�׋�#u������K�	�4��N��">\���+׀��3�~��um��\��hC�QD�t�t��`c��Z��#�LnC�:6P��Ԣ~z���r*g���-�M�KJr[�Y/�d�D.*:9�x%.)GH��DC���ZdK+�l��J!�'�*�N7\���)�4̌g�� TT�v����Z�^�@0Z	 ��#^]Zqs(��k�d��[�3��.T|u�p���̡�8��~�l+�M��� .����Y�����1 �?C�*qk�1`TD�&!�2h��3��֢��z9��Zr�a�[��h"�V�[-��~q��Q`�
�Y�\R2�������Y��{�D�G�x���u������r���ߣ�l�7�0;�1��  @�w�s��I{�%����[�_@��ov|���E���Z̲%)��ز�9'������-R�q2�p�!G�{._���M_߉��b/����<�8l��H�t�MD�h�uU1[�c
rBֈ:wz1��vs���6�RM�o��\�d�n�,㰺�G��]�mr�Z �_H�L2�i��֢i�Wh㦦>#`��\����4�#nĲ���O�a��`%����J��pf����kpz5$1��w\�8Or�)'^���L�bM�$�0#8�K�ٵ���1F���ǴK����8����+�6�ոB9��4K�m�_�e�TWx�{~_%f�pU��P;�g@����#���Ku1}�_�WBoצ����Lp6Q<mr G���;�9�8q�$��^�{���Q�٤/v�J���B_�B��s"��c/��D�q'��r��KhT�S����o	��O) ��]FpV������ �f�L��Q�z����}y�'��ޥ:E���O�}8Pb�VSN�J�� �ȵ@k{_]��,�������k�:Ǧ�2"P�	"�w%i�4��w��&� W�s��vR�˗�8vw�`M���������)�O�O�#�U��a#��Z���F	������'nW�q>K- �i��[5��] O���>(\��R��C�6�A6�
��uG:��^t���_�[ou�	S>�K��F!�����:K!��� �i�|
�1}vX��Q9�q����O*�R�g�����R�1猰]�s<�H��n����t��<�I���� e�
�q�@Hx_�M$��l�2=hu���P�O�jEnJ�:羱ܓ��3S�^e��X��X>��gX���XO<�z��;�:;�flY<��X����o �T�����Ԟ�$_������nE��;�j'�p79�:6L��D1A��fx�AD���ːEB�>f��!�؟�T&'f���K�i&ȴcl��-T6�g�mXP(��}�;���@�:��Ux�N՞�ؤT;��~��I f���ۀc���<�ƢF����w�Z&y3��@�K�=5}~��R���0�0�,���Q���|��M=�����η����M���Y5�9�=�Ł��C�iu"���ˍ����qد�N�����ˋv��D�Mr8;A�P։-�g!R��+���f�X���K�:N'��S���7�<J�n�0i�}\β5Z�K(��m�yl����y�"=A��.k��=?�|�<5*^^ei�1��pefO��k^���q�����VRx��O�2��k�Xw:���D�J�~��S6��e���^3�d���J�d�P@^�C�\�����o��'
U?�z�#֌fa��R���*�` ;I �a��{_��9V�#��1u���1�8�ӂS��W�N���%dF.�L���qWb�yd�w�.p}H��^'����m�?o��8)�����'����Y�ן2%>��<?:��4���7�9/.��>zD���;[{93�D����ădj�	�ռnmaP��2���ڮK��Ű����X��z[�|�h'D2ֱ@ 渿�W}�1x����w����j��$f�!�t��Ce��Z��T�Z� ���g���޹�N��sn����y��R�_��bD�ߨ�?��Nr��/UOH�
Vn�]����S��'tB"i��y�p�j`�����P�����)��jSg��|���O­,'�[x0����Ͼr���T��Q�	��3���4��|�W>3�EP=���ʝ�|'�n��ME31�-+R��?*����nuz�=u�N��K��Z2%6�Tb^��lw03��E�O�1r����V3~�+��
�P{Ş�~�DM�ҎY��!�ج"e�G������hb���s�}&`%�K�>�����󣯶��:�-%�]������]ޔ���)�>�:[cN��EM`P�J? r�C��v��O���Mp�Zظ��ȓh9�$���ʌ�-.���e%�Ӧo	\U��bV����%���D�Bד��( �T~Ȼ�n{u������ϒ�B1G�&B��S
�-'(�-@��̂M(�#,�>��)}K<���:d��o����²Eǘ���Y[X'<�?!=ǌ���M��Ec����c=���j�\��ڟ���e�&+2|�>X��)�Zw�V�S��%��ڵ�0����K���Q�^P�BA�lMZ����~%׹��,)��ߊ"B�x�X�y!	/jߕ5���*Y�^��WA�ڗ��(b���!}O=���a���w�B~�V�_�lg��P�>^6�n�	V�~)�_��h��4Wpʶ�_g��ҷ�Tq��z�J��-���'ӑn�H�3���#.mw?@tE����iSIm��|�k��GG=l���;W�NB��,*�2�t�-w�#A&,+���g�{o]-��^}��7̘��bm����`��<tA�-Ⱦ~D�|�
<X�#�x(�K��i��` �3c�g#������l��yV@�-���������^~�2��	3��� Q.�z����w�Ã���"y�jj������V�;Z�]���L��%"���k.�n<���uڿ�R'�&|�6a��S�+^��r2��fJ�>M��p2o�o���bN��6�c�:,&��f����ҝ���F�J �k� R��M)X35W/�h�E�HE�k_q��Ւ�B�-V�_��������&�O���$, M�ޭi(�+��d� ������ ����&�`�;7>R��xp��o�_tyq�u��5V�lE��@Ո����v}x3�)�:g�MK��&7�B�V���%8�fy��"	G*_gӹь�^�;�L3C�:��+48�ϘdZa~o�L=y��e�\��m� �<*&�kJ~��88��&:-<��ٶ;�[�-J���&�l$��)B��7f�E����z�'+)6���$ZC�$���y,Jߒ57�6#8���#��M�u���g Gd�6n.���99<��FW�=�-��
?�����pL�.E�?�� ��t�Nt�>�^\�sԙ]�.ܤ��.�66_�Kѹ-��N���a��
�C�|�SՐ����1�~�����P\� ��I�6븾�)�]q��P�EpZ})全>_�O|����c\~r��5�1	�p��2�_V���m�+�Κ�DM��}IC�sX6�=JP�XS���0I�����ݤ?�>hZHi|PJ��@FUJ�)��z��`���;�g�1��Y�G4���&@;5ѹ&��|At�:7|w�c���8J>Le�ϣ)Ŝ�{N�W�$��-���v�@�QZ�.B��0���ܥ�֯�Gz��A��U
H_���	���_o7ի�νV�Oe[�T1������)i.���a/��<?��\jt���Kf]qG��B<%��P�.0O�<�P��;x�M�
#�dX�g��bO�f����H;kz�ĝ�����*y�����]B�^��W�0����"ʄ���"R�������Ķ�A��o��)��\)��ü<��[��{)��I�x����?D�}�\q�X�hs��B�5׽R���;����V�m9X}v����n���k*��]B4�~Z�o-@�B䊵�3n�d�ݎ�}~�
�/�E4��	��Y��~��s���<�ƪ;�C�m쨭��gX*-v¾L\���<K[G��bƣ��r��n�I�Q�ن��NHwF���K�oΔ�M�Q,Q�8��
�&[bN#b�Ix��V�3��)0�1v�62���.��O��9t��j@�,��qY�A2%{��A��Im+I��T5�;%�҃{�ϜN��*�H��3R���0�����y.!����������:i�up�)�'�f&Ӵ��?��h��;�̹Z�S@8<5��C�x�'6o�V!QN�rX�� �Ꮉwd�*�u���zf�A����m�U�9����e���:z+�6�|���P�>g���-�̤F,�k~��XPs(Ɏ���f�z�	A��˛,�72X�C�X*�u-?\���<��x��f��X�sKx��8�<������0�u0\��{��}�Y�'5Ų
ۥ�;��[����w��g�L84l�T���S�h�Y��n�����#������z�-"F��C��
r�d��G{ʩ�M�)ӏE���Yt?�3�~��Toż���-qA�w}�.��L���B|o���&�f�F� /��,�3�n�Q-� ��X�t\����C?Ii1�O~���9SY_����+��V.��B�%���T��5ƕlk]׈B��g��"֖���1ѥ����FW�<�g��>2�(�ǹ'���k�o�H*oe�ֿ>Q����2��5�F�W�QH.�D�Q�}=�U�*�8���)<.��q��ߥ%�&��-l�i����2u�����0>�U(ݥm �W'������̿���ӿ�U�����v�Ws�p���!Ϙ��q�ub|����W?;xK��9��,���d��