XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��15_���&�4Wka�Z_<���jo
�����~��4َt����\�i�JL|�]]˄P�����q�V���B|�A�������	y�Q�ڄK��8������V)�g�y찦�H�g���j��(�ghp�w�Ck��<*�m,���5a�j�k:���Q�!HT��u�_V��0L&�W;��4�����m�\��?��n����0��7��sK؃f�=o,�2�^=-�瞔taf��8gN���7��]� f�0+���v�7�� �7�V]a<���J3,d��B<=ߕi���RcY5�L��i�U��1��	�d��ѿ�R�CbI���M-C�2$YY쾑��I\sz0*���cT�k�g�ͣ]�C�q2��h-NH�MI_�Y�w�ف>}\���_�]:�RC%�wA���e�M��F2����F�2(�3,���ƜE�L��Ĝc�Ʈ/�sM�v���Z��#Z��C��o,Y�����*^�����C>����>��k���f�z�#����1GZ����?Bڥ{�������Z= vB��!Uf��j������C���ђ9�(.[������&�0+G���� �ON�dO��.R�Y���cd#N�0fǵ���Y��/;*�V)���BN�9u�`���D�a ��:��g�WwM�b,�1��ۗ>�r���fiI\�d��`@*��"m��m��{ ��5��3:����P��.�[���՗k��:{���ݺ�Lnu-�P�|`6��u|�_|ڋư�b^+ۏ��XlxVHYEB    17b2     880<H�eq��`b��J��q���G�U��9�Fk���kJ����]�W�pf�EϪޞR��\FӬ�8=�RV�^El[[�s�M��Į�l������b+lL���!H�Ho�.�n	��=�a|��Xۉb>�/���W���PS��	�fO.u��1R|�3K![�Zw`��۳���'��J��@Y8�1o��5�ƿI��aAnC�0�_O�h`���gH�)�S��'��@��a�[�W<Ik���y>��s��cw
��t{5���}����r��^ߊ�MN��hy@��`E�[UB��;�G�+F���n;�^��Q8lX�l���Jj�/ʟ�c����)9���X��(?���<������3��duPvx�щ�Fq���9yW�?!o�B�Y����N�ƙ_�*E	2��1+Q�tUf��-x���_E`Wh�4#lc�����1��$�䒺��
6�=��?Q�D���W�Y�0���e�Q7B]��+}��J	͒hY�>b�7uۓ��Ȏ�+�g�\���
+"J"�2��?�Z̄�;��w"�� (�lU���^9F�~�z��@s؍���P�ذ���9P��Fʯv�A_YV��K���M��9f!�2���>������,�@67�P��;cK4&Q�V�J��4h�d8���6)�c,E���Y?h���<�cٝ���x�<t�GD~XB�? G��̦♅N4��Ϳ��u$��D�� 9O�8����o�*Z���D*��?YŐW�U�RK�S�,&Ϫ|�8@*n�����A��}�
���V����۞�F�U�f<�ATk���5�Tb��������Zd]�{p��K~qw�L��me#��d�G�66[?�_m!wiF�i��`E�F6�E�)�R�@g�a�A�rdꂩ�vD�wбnCJ�g^4ӗ?��s)��{(.[L�*ڵ�V�ek6��#�������@�7�Z�V��9�V�g$@�����:)��$%�3�͜�SI�-�� �����W������0jb CD'#���U�x8�����@�67+�$a��d�*}K�{^��6��`7���w4��._
�g�"k�uіPn^�N5��W9;�V�Qo+qڻ8ԲKN����0%F}E{�ĳ�F)���([7����e/��M@��چ[e�����lLf2>8�j� ze�RX��~�����u�&�nr%��w	5��z� &�&�������H�OU�X��DpL��%P#Ӷ������
Xp��q��)
X�o��M����:�� �M�A��;u�jXw�!_�ƟF�1�_uvCʆjJ��x�Hn(�iY�Y#�g�3?cg�����ZY$7uDD�xj���� o����3�>ҟW��e�E��a��*� �Y_��B�Q�[F9�K�Ok��s=7��%�1��F������3!�ԗ��'Ң��w��W�u�2��2��˶�bZC�\��>_��Q5zI�*jBK�p紤���/:�kx����� ����+ �� Á��Pi�ڮbOs��]�΃G"���I�	l���Y9��b�s>�/tF���xv�)���W���dk�@�Y��� (�юݱ?Pb�E�1���ȸQ�)r/(�2|{�Nr8�L�t���v�%�P��č]�:�������Ǥұih�C"��w�j�b
�u�8��������w2<��eQ�;�����eM"#[�w��~�̞����kh).����j�)�r! �XH}Ni�A1�F; �bp�$����@v�,I*�̡�}Q��?��,V�~SC�Rx =��d��~}��HIEx�v]�n�$���O�u�V�?ߗx����c��P:2s�����)_��Q�E����Нd1Z�0����GQ��]���x\����q���N�x���h�a�%Nt�/��Ί��H���fhR�ɬ��qƁ�YmS�q���m��l�9����h&cc"�j(k�z1ms�� m}�M�=~B|��)�;�oZ���э���A�y�|ôoU�?��l7�lCw�DT֯�ZR����>ڈ�����8�jJ�n���<m45�#=^/f������_:)D��I_������ij�q��.I3Վ�:�^�9C��|E�:�l�
