XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������Р�'�*F����¹L��(!E &l���IK����K�}%l_��6F�%[s/F�Kw_2H!I�i��݃�X��WԏXPu
H�k�T?� �����!��	l���+�V� �Q�9��*��)t�bsV��"+T�@�ނ�r����]< �%/�Ϋ�|G^bO�5K�RVÝ�Yq�`.��jM��� 
ёf֩�$��`/9zU���T-���X��"��d�Ƞ��&`"B�@ͥy��
���r=�k%^�b�`�pw�_s襖����&�����9�����y�
b����ϱ�k��R%P��t���Eh�YJH>��g	������ߕ��&+B����s�7�G�`|�=oD�H�|��I㖃\����ZB�}f�iԠx���<M�,�?�%���^�]���_Df#3D@K|?od�֡�M(��
��
t:>�,w�3`��ZJ�C��Fq��C@6���v5�[���j���=��;����xF��1P�a{d0礴�O�ߙX�*��i���9*�QSZtȁm�ca92�|�&K&~�$fsm��p��Va;ˠe
99P+��i��udm��<,���-*�wuj�^�����14���;��3w~�J���7����V-�N{��:b��G;AR�I1c���P��k
W����a ���J��oeEmYXJ�L%��JR��������>�����f�����쾤F ����{���3�dử�A�0��׮Ǜ���]�����S5XlxVHYEB    15bf     890W}ú'k���M�w�;�a��9���I��s:Jʫ�b�4����
E�c(�&.G\�y�7��a�|w��[n�p�N10Y�coSmn��ֵ�8v���9[�����Z�B�$����v
]�� zK�A	�������R�f�g��G��ȩ��! j�7�?^3�_z���E�vJG+�M�6~m�9n>m?Y�� ���Hӈ�N|^&~Eߙ�]݋��!\�<n,�r|�7��j��Z��?D��-T$��<(��5[R�S�ef�]��Ye�[KS���
��v'uX�/;�_������*\�*d�)hT�ґ��G�+�rؙ��b��jԨX1k���#��N2�|/���Ld�D��2�tn�~�/~���t�>dM!�%R���w7�(!7C�C�s�_X](�PG���0���҆u��{�q���D���-�q."0v2��H�b���+�2u��U�c_1�ɂ��SV��{�\!��o06Tje��p�P��ʓ��[{����X��@tg�l$&�j:��#�ľ��Хn��²�G���o@�[�=��U��������l�M8�jN�>��љ�GMA��/v��c���o��.���5'=h��IPе��W$x��S)|��x>ju��6�b�E3�ؐ��/���N@�[8��(fdn�= ^�1�A��)�!AV�=f�Κ�8���{9g�0;��gC��N��8�<�%�j�	��^S����l*q�}�ʔ$>�+��Ti,�̨44T�(�O�3�LM�'�V�ظ�0�p,�.����w̦�bm�^�c\���]����������Hu�%U�����!2�'ꛈ�2e�b�j����p�X>��+�l���"Y���c�ڢ���@�%]��}�@�W1���9�\��gǶ����?��\��?�h{h�o;f�xJ�+��25�s��p1��6#G-���jP������#�{R���v��<��5_[HX3&�7��RV�6�(��9xö)d�[�A�̝&=B�r�tO�A�ߧw�`����i���))��ǀ�6��	��6����3a�ED��62-\	�e���t�ƛ�Z]�@ &b�f�}��r0C��!���F!��\Xp���G��d�WzM�}���~?-K���O�Bz���t�[=��Xʞ)>�\X��b����J��^ "_$S�kR��]�~� ����W:6�lfz��:F��6�M(�W��ҼK�l
t���[�𶴷�~�A�5�8�:F�.�3�H.��>H�+D�N����� *M��v[�h�lܕ�����	�~���o�B����M�_i�@��s�Ǟhx	�� Z�� �
��;�{֬��!�{�T���-��G�|K�0��j� #K��rV�2V)��9{sW
g����Z��]� വ�hz߆�����Z��;"�'k./ޔ(z�ܬ�K�r-FN�6�gx��
U��g��󭟞p#�p��'r��C���A�\M�h��� �����Q�g�#�Ѵ\�Y���h��mle#3��C�Q��<9�0���W���ȳ}Ve3��)�a�:�9oM�F9��[��Xrn��h�4$5М{�V��" ���Z�9��)�ɖ���D�_����)��@��z�!��7|:,
JBWE[JF�`Lq��-��IfQ�4�W���wl!ùKP�h>�9�J�N,{����^�t�����'�h
ZϨk~�׌g)�
�������b[�.=��z��6'�:����##�ʌ����GH_���{�H�{�pKv5B�3G��7��z�9p�f� K�ީ\z���}�{�F��n  �m��$�����}bbAU���o�O 2̩d���Fڭ�Y>�����S>��e��[�=/��x���	�p�cRT �if��~ ���(�!'q��>?�*,9��"NwO̘w��G����UG���3C�s�������CZ\��}�b��f'Ѡ��Ԟ�Fl}��	`�SF����A�H}H�6�'O��y���/;f��4�2���(��MP�̳1z��J��J
V��~��e|ԟ� 93�g�ґǮ����.��]]m�V$�N�i��F��ñ�č��\�'��T�7k�fl)<�<�ڡ�m��4& �#QǗ<��b��6Y��jgޞ �(�1D�@ر��@?�