XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��}Z�[��3>־:G���+��V�\֢����Y+�ޜ�*���숫"��#�ؽ�[��4�6�5�}���R��o;���H���MZzp�'�G�������{Kuu+�+�~��)ŏ�u=/�P��$�@�x������ژh���!�!�Ò�N������Q����>�ę�6f֨�EAYW�����/f:s����iAҍ��n�e0$U���:��>�+��mB�pu��:�o�5�"���z<i=E$��:�@ ���C�(ӆ-P���&`\�,r}1U�rέ�IA���X�R��:���{���8B+��T��{-1%n?�G�s�wÌ+~AHW����`yg���l��y]��=�j��TZҊ��T�Ͱ|aQ�f�3ށ�}�*G�i�D+�A�ɤ�,>�Q: $q�2uL�0�K�P���АI����&��R;�À����P�K�)7�y���Ѹ��A�+v�p����3�N��3���]�=K��� ��d�r��/��<:8ҵ��zV��o'��I�awrs�k�����8RD	��$Lf]g}p]�)����,U�q�����C�5O�zzw�2t3�8����b���Lk��qC|l\�xTsxeOD�W�w�nt�q1���>l,�]MZ�SY=IA�w���U`��R��<*haM� C�?Q.Ҝ�c!�Wl���	챂�:]�����9��H�T%��3r�VR<�-�7����XC�ê,y��g�tHR~u�dE1X��;91Q��j�X'��!'�XlxVHYEB    3e93    10b0>��ud�(+��GV��� d�v��I�쿤${A�pJ��'n �y9H4 ь�(�8z��\D1z�az"2ݛ�zȪ�l*Ӑ��G�ԋ�t�@MLu�F�(ɢ���Ls��z-T���T�hP�/tT8�n]�oPF3�וR�g�~�*@�营�����p�3\�s.��^ꓝts��P/y �n�n�&צ�fU!�
iD�����Є��XV�� ���5�K���!R��C�x��Y!���(����؁��o!�l꠭��0� �C��\�j�ZV��y���v��#� �ڮ��E���F��HMra�`7����˵�{�, +ݡ m�8@� �����?�X~#��%�n<���ػ� M���ƫS�`Q�K;�M���!5׼.��懻__�\�V�T�&0;D�P��ǉ�S6V��������|逊�~�
d�CY�����[�bG�}u���B(q����[�1(�����)�;�7��#�iמ[�>�����HP-i�c_0h�_���Ȋ��k���6�+颅>���>��m!A�B��@T�

�_Es�_���������W�9e��,�^��;��h�`�����GЖ��Q�^K�f�C�3҈��fs������Y�3Ӎ�7`��S��D+�:�U�;��<�2غ�=��Ϝ����ٝ���7=�����p�s`�Dg�*�3�U8a�$��w������mi�n�`�s*a�Yb��N<�+g��v(Sf$5@�r~ɏ���e6��x��!��Q9C:�:���_q�L�%E�8Cd!-�[nɝ���#S��?u�%l("�g𿮛[	v��tx��|
o$�׈VֹVĿAI���z:"��3/�slQ��/���c���RT���QBdz{ }��J;f����5�먑�s��K��q������c��r# -�N���oʗ��|_���G�DA����c���j��Dw��3��l͇�e�P�D�U^?6���3.�.|R��q�)vuS�����}qW��� iر f	z �1h-��2�(��($���\�����V4V�E�p�%w}��.���k�cG%��W���.��C�6s��a���n�Py�s�*l"�D���N0TS.Kq�=��|\}�ݵd-�?���r������r+`8t�C��
�Mih/����s%R���=���()YQ,̤5�e��T���4�:���M��q��ۥ�m��vl�}������Am�DW&�'xb^��$�<YA���L��}ެJ"+��\U�PA9��	�<;:�^�?���H��4�3��j5�{'���lLk�t�h�il����㵌�U�U]H�_b�)!Ԫ޹}���\�|;��3��l���������LXq����f��hV�7�d\	�u��bX�>��߁���}V��Qr$:��s�mw���%�ݡ3u/�9l`�O<��f��W,
����>��\�SYӕ)��˻ݴ�.޽W�[�p�_�r��{3�u����������@�����u&H�t��yq2�l�;^��{~���//��"��i��YOVnv���KIj�˻����(|�ƶ���nT܏�7B�5�)�W����?��^x�	���3�F6h����n0<�R��/���H�f�-L��yTF��RG��N��H����ն'�ݑd�uk[�7R�)�յt���?�'�W��ܯS�,�I�=�_$��\E�mF�:>� 斢�yP���h��h/4w��D���{i9�ԍ����]�x��q6�FI���i)�z�IZj�[���n =84�;�;����H�q�:���Ò�@�mg��?�.Ұ��3�r���6�i�[�eA?�����!���јH�ay9��N�}W���txap�YT��1��v?�|do1r����ݜ�Cc'��zP&�(|_�n$>�7;�ţ=��.y�G���}(u� +��/����n�]J��"�\t�_E0[o���W���,&b��-�j�@(њ��J���~���^�	���Iab=wK��|m���j;=S�� �G���5S	��,3$	�o^�O�7N��4�ϟ� �ls��'���I�=>!��Ya�0n��?9���V���(��m��U��f��D_'��AV?�5x�eȻ�&aSM�V:���I7�/�Q��>Pex;PE���5�FFX�)��'F��b���k«H�P��^$~G�m�+v�U��]��ž��k�ݟ�2{z��ҥ�����p�c]���x3�L`��]���(�އ���&[qi�_A�KG#ðk�������usEyW6�R�6ȱ���܂F��/G��Y?�-G'���Y��/�˗�H��DZ��%9k��7�}%�X���\}�eg騈�b��v���D�M�6+I�1ğ�T?[S��$�`�@~P�3�=8d�/��cF뒬�tS�ۮ���c
��+O������+(��]�����݉@$��#��`���Ȱ�s��:��,�����r�M��Զ�Ϛ��ȫ��w�) �%r�d^R�)0:�OE%@��t�Z��q�K=���BO����4���(�i���+K�&J��c��d�Y�i]%���"�I�P�[oO����q�x'�G�-+�38-D�
�zh3"Z�,w�k�7g�f%��^���-�W ��h�����P�+W��1�Cb�ק,�9n~`��|��YV[g-7�vx�f�2u/̚ߟ��P��I~��N�{��Kr�(TG��rނ[8�,BH1��"�'�1#�$9�׸���Z<�L��H5�/�|eȈ6�I���A��HN*�<(l��*�ri>k�z��_��K�;�q�n�����~��I�J� �]���l��۵yܷ ǝ~��ݰ�4��{`	 W�� ؗ.o5:�UN�Ķ���)�� ��<��8���[N��h��Y�'��?��� ��ﯝVC*s�u�u.?iS� ���=�K�!�H4�%�1���	���D���?�G4�ۦ�r�M(����.�S]g!h����@�����O�ׇ5+C��} p�&�9�S��K+�)�t��n/�2������A+�d����2 1:�'�8�gwNf��X�u�Ka��H�|���1��]c�>��A�G�?pۄ��~��$,�m�Jj���̀C2���`�Ď��ާa�Y���~?�$��RE�t꿮�}`Rx�[Y����D�B	=%Ǝ�3a}����͒��b���~�
�n�sip�]>Mb6	��VL��'C�G��f1s�Cc��~Eu}ذ��y��ꕟ�B��w�����Σ���)����B;�5�wm#����l�<�m>����z6>��ŠA��gL�==}}��m=%���Z�[���Rٞŀ��E�+��5%6!�Ω�x���]���K8�h�֢h�d]i^�����f�k{��7`E���n��J�c��Oq�pv��?��mA���2	R�ϑ�jV��ת������L����w����ޡE���,�"�s�`^�*�TF���txDTe��k�'��c��6��2��#�G/Z���Bע�u���al
����*��*���S�H�6��_��
{��qiZ�1�.��[���Ey���蒤��36����ۿM+�hRC U%7_���@�[�����z�JGP�s��]���p�d(�{�^P�O� nl9���m�H��:X��e�%=�&	��g9�47�y�Z�\�XN�x����S-������@���B��-2�M�|]-����3Mxz~�PJz,g'_�5]U ����d>]������2��_u�w]���7 �-XB�O�eë��H��&Cn%Pz2�Ǥc��+_`�e�BF5�y-Ӻ��y{��{<�t5��T߫�]c�twͱa�9�S�L���e��t=���0ꚑ>�OU��b0GR�۪x+~���]�fOd$���y����R���W�i,g�H���c85(+��R�e�u�9�����6x: � �X����vY-�v�����?�y&bl���"��њ�*�wL�Sfd,;Lt�g���n��C;`m��C�Ge.7��c�yn��{�Y�m�jE���͞m�n|kVW�V��� ��˥k�oG��)�a,1+x+����c�ژUQ�m�R>�z��� Q$I])"�Ǥ��i�[5Mu��>�Zz[,����z��DZz