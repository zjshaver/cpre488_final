XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���+���=�^
��D��ua�e�Ů ��|���b	��m�3x�ed슖i�@4���Y���_n8�O�z$|��-��{��c��Hm�x�����	��vE|q���/b������r�n
X�Ux��D._��+�Z8��bUR����@p��8��Ґ����O��ZLw�3,��,�W+-�.�F�\�b����}*�?k�8��k^A����mx>�ZZ���I�+^����4N��+����bГ�뗑؜��� ����~��@�3|��t�A��+N����<�h��Mu��ߥ.�@��|�:ml��
�U�ͯ{�1D�E�JLDJz�]�.`��@�S�dA�A���|�me�M`dnr��p����&���PY o�����'����_Q?���?u,�V͘x�C3ɴ���!���y���{��y/|�|������l�� �͘���VL)���̤�9��a�-�sx��W�����N����BH���Ծ7�88���F�G�/��w̫@�1�bsӥ��Aj��ϫc����T��HW8�RC���MDyB.O�v��H���om���]�r�^���0P���$lB\�ܕ%ͻ�� �6���k�"�
�w�7���K��4Jj��˥�4����d�E�D�'��m�Zg:}:e�N;r��1@�8�Dܳ��pD娠���e�q�P�m:}K����t��&�V[Jgq��E}�� �X�qXlxVHYEB    2b39     b10x�`�7�x��og�1ȗS�oa4�`���p��Ut�p24f3q)W��#���4׵'YV�H\�L�3�n�E�L?8r��`�o}
��i�2�ҍ����P!�ߠ�f3.�+�yC�,��`��2�&�,d�'�&�h^�!>���g/�����I�$��1�[��슘9P_�?�n>�+��Zx�����7�"W3q�������ʓ9.�P�
�[�@'��kT�7}�����~Z]ē�b�����&O����~%�í'�(���<���]��bɼ�֝'�5����*=�v*_ٍ���ߡ�Vc^?���gЫ��b��qO�����(�����)l	}�r�.c
�E&�V�x܋p��	!�����s]؋qSN�jB��9k����m�Po�3����<�2��_{f�S���3�)F��<t���z�����Ve��y8��wlW�/^5�P��ψ�g����ȫh��R�9��Uu�������/--�,�D�T��W�h�\(��YNd�ˡ&e�)���{R�#�Y��:�̂x� ����g�.tY�?��Ю۬�o�6wv_'	�S'vg[�k,����>�P�ʌf�3o�my�?.b�C~U�;��M{��,���.���U|r���nZ����ɍ��j�|_l��LRX	z����8�������J+��gh�|{���C����P߇O���گQ�D./\�XK�L0T�$�ƹ(徯�2��a�V��,f9�xA��S{���Rpc ��46�Y#�f�"�wL��ҶK����k4��j2���1����?t��<}_jL�L���� :j@�\�x$������/v���NY��mV?�P��pA��9~��T�9���<��IZ9;�E���{c���;��㹖�Ă�9�v�/^�H��O�	f�f�<��Ak�I2���L��17�KIڷ�!��4�H�YFH�>��5;��V��E+J��>N�!]���aU���p�,���Sq,W.I�=�)]J��%sz��c��>n��ѐ2�~�{~�c[[����5�l���{&�����M?���~b���"C�Z����3��K9�S|�.������v�aߚ8�BCr �������0[ic\Gaq�`�'�{�$%|��7w,���V>Mq���M.-r3.ߍ̿j��./��W��O�� �xn����T�v������Kv�$L�6�$CM��p;�E��i�I<�-���+�&-:.3�.̳�2��ΧQ�n8��=��eD��]+����f�ι��@�{;i��x���>�l����넡Í0�&I)���\������ּ�~TS<gS�>��~8�>�3��n�H���t��b��� ���:\e�J"�����y�8�8�a���9%������ٹ��1m��K��t!���틈�Ky��	8'�����l�\5�>2����SYS�m39Lڔ�nѧ>����Q�ֿ���fp����M�[\$��B^o���;TX)!N\���&n��8~����}�̙��kE�C+8��e�\&JE��U�д�G㖛��pA��K�!�l�Fm���>+N�}
o��ϻ���-03���$���'�DlF{�*��E�v,p]������:�dH;\�w���FW���L�"�.�_��+�n��<�M�x�,K[y�k���A����o%A��0�q��p�Ng�`W��	$���#��y����.W�&���í>�,`&à�)��Q}�C�w��K�������MQ��,%������G+�Ѣ�rV�%ʱ+	�CfO�nV�p��b!��ڰt0��vQJc���-&�q~ۄ�]�;�A�x+�a�w������0���n:�K�3�<�5!�W�w?y$�n��<�J��q���"�3N�ܹ]	�d��٭�s�Nj�A�l@���A�c��7.`�q��F��J��$��l�^=�<�L[���cr�ɪȺ8���U,ރS����O��գ��{�Q�|�^�Ǳ����3�h(��ƪ������*!x�k0�3���j���#v��ֶ̨=�C�ǅ�C�Z�ӳ���i��@8���^.�o�
��p��ev�v���j��K`�Mo�d-�FW�t�1�*�}����&@�t��k��
�p�kV�k�ڑ2[�7�8�P�*�s@°�����kГS����X<2�|�q�@Eg�(p�8���^���-H�L��wjGR7fTH�ؗ��><]�!k4H@�cLg��aU�`�5���m��kŴ|^���17GG)������DZ��(�ed*x�BHQ4���:{,v�L��Ѷ��f��m����9�6V���������h0Q�.�� J����/M����j������I�6��l�j(�4�KN�λ�Q�b��ɡ5�#���@�1E�1XP��^Ҷ�����&�4���
vl�m��M��\�2U��K��@ui,�
���!ٌ� 5�:y�����t����+`����K�yэ!2A���YGe	��C-��6�)G���O��E��^�#�g�x�H��i�A/�?�O����J9��$��ݝ�T�;��dxԊ�Or2u�٥Ԥf9~h���mJ� :8п ������ƭp�� Y�`�M�V]�Xy!Ǌ�{>f.���>���3��Ll�9�8O#B�{t�( ��C�(�����@]��<Lj&�'�{pY����ѹ赦>�hr�k��M:궰h��2��qY3�`~�f���b�0>k65��n��rM���{� �n�~�M�	���e�3�