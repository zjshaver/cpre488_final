XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��		��J@[�O1���jLs�=��TLAT��j��w�{�l(㨓���d׵���o��;��K�)��̚�W�3 J!����#3�<W��N�Y�i���Q6H'�J�q���-L�
�Ⱦ�8�F���iyGi�D��.x��x��8v\�������=lߙ�`Ap�Bj{C'�C�ƒ�5���(�Ŀ�2���aX���{�u���k��#C8�`𶵨S1�+!(1�א��WA�xp����E��x��j�K[WR׆@]uW�Ӈ ��!�� ������@�_;F����0q4i�M���:�U-ɔn�����04l�"�]�~Uί�,7=���}:�f$�;���-������ЭO��P�R��/(g�E��p��X׮�A�j�����<7?s�Ç�"�)�b��$�������%:�2ʂ
�4z0g���'�R�� ���䅧1�"�jL�y��a\����)W�5��AW�1u4 �,~N�{�O���>v���@�`*%������9�[�Uc�}2�Y�q"P��͊[4Ŵ��ɚ��a�(�f��Hw`@{Ò�L�aVs��p��'v�W\I0e-�4��9����s�� x�M��Lۦ�6=���3����Wv��7s��ܸ$!ݖ�-���$�`*� Hw�k��#u�?�3���D�htɂͬ�{������X��)\p��Ui��+Mg�c>L�X�� `���i�;���t�v]�H秞�(8�c}�(`H�܄��hG��?c�ء �{�rO�8���3+?/�XlxVHYEB    3b09     f80[Ҽ��AMIb'||�NWZ��[�UЍ{��Iib^�.�2f�;��]���?�`����!��«oiY��C�":���;|N�%k������3�7�ed����e�!#�9�(g��6�{p��pgG�)����2����ZC��VYC9pQ8/��E!��Я;���pko=vg�m���ܓu�aã��P����~I.�������`��oz�P�BB�u�����<Vv&w��ۻ��ԩL)<����׷��v�&A�w?��,���|�����Cp&ˋo��/P�<�ʤ��a����G�>Sz�z*S�	:x���I���w���s'b::IP|�aW��n�Ϯt֋t��zN$�se�v�,c�����Q=�~�
2��,���p)U���({��1%���>_�j�/֏�p�eZƟ]�w�Ud8���$��
I��kЄ\����e���r8���q���d�jf|���i�m)�9z�MѸS��NΒ[��o��T�1��Q7�'f6�}*b�'N*<y	�[�+�z{�	�R�ֆI��&���F��:���Qq0j�1l�1��8�F�邚}Gx��M��m�b^��hg��$h�J��3��7"��T}�À�PW�:��&�2�8d/mB�Z6o޽Öq�Yu��;�����+�����S�5�N@�l��' �#d�U,ɶ��[|���8����e($�/a�W�q�����ܶI������gJ۰$�M�������vlU��O� ԡg�%�����r��y-6�k�/)����/�����<�^�+Y4�R�Y�&Q�!��8���r@����ֳm�A�2%E"���Mt$�t��W��l����-7c��A(��S,��=�G&���"ڴ��h���So��R���p\�ᢞ:N���@r2�D�Gj���P;����5^.)>2���C���3�m(B�ł�CXB�k������&�b�U{t��IgP,��4NU�>T��v�� �N��:O5�&�?�?(�xoLp�S(yԵj�"x��u���a�a����d�7���Z7�Kc��'ا�&����+DifBoY�X�C����M��Cc�o�!��E���wRH��r��I3.��J1�؉xj�[�A-�QtW��+��>X+�~U�S��~���	%MK�K�de3+�{��U�����%��z��뫭5����`�����Ȫ{x��[��s�,� %��cxAF:��;���w��-���b�;gCS�'0�8��Hu��n�j�3Oa�	nk{�2��VOR��:i]���K��i�(#�����V0�+-ϼ\s����V����G{��li
�F$?�î�R+��'��A�;�pq��1�5Q�uKL�gU7T��֔܄�*m� ���+4ݩA��sOW�`�4��0Z�wV�����*��.�s)L�3 nv�p�0r�o4)�ƞ��zoQX�­�?�p.��L�������+�NF�ʣ�s�3D0�Ja�KC���I��V؁/�����ÎUo}�)Y���b�@~r���C���ױ%��9j��F yy^���Z��x�1:B1��S/>R.
�|��B�ܶ*
�uBժ�ލ��Q�79 ֙J3��0r�lcz�3Gtz�����.����V��"���}/�}`�Ե~��1���&�S���X�.��1�mp(����ߺz�g���X�aބR� ��hY �l4D[YRz��l<�*�e�������ʫh����Gd���k�:�U{��V:�e��<iNDS���v4F%�ɂ�JD��`(���0�N�7�=�mr���n\=%�;3� ��5gζ���?HͿ�p���Y�a�u5��H��uW%�_���#��ػ���{���Xo�?wW�~5�[��)��j��B�p�fb{$j�su��:g�H��He 1�m�c���*�Od��ɉ���#�n�4!�\�����H�'#����)ћ�
��¼
����$'}�{a��W1�ԋ�j����{>�UV1$\���s)�8,��3��f���$t�.��0��ӕ�~g\���_��s���d�<�;u�� ��h[u��~�e/�Ĩ��R֙�LF�n�<]�! �*�3�F�Y{(p���)>w�

č��*��W���8a%ُ4�?<�J]�8ݐ�A����d�7�o�z������h��#��ړ����ړ1�33>���7�J��p
;j�z���?�J[d?��\]0$I� ���"M*~0�&��B���ӑ��Iʫ}��� g�L�P��"��9���AM�����,0Y�x|��4^�f��pV@	��r��H�y\\ұ����&Ӆ�3�Y	�]�S[1�&�്��N��X�ʱ���$?�bB�|�֝;jޝ�O��S3X�EwAe��X z8bG�E7 ��#�d�?��FS�(�J��=E�,WF�#1k��Q�w6�'�T�hW�$��#;@p�����#�/��Q0߁�&H�g#ρ���y��̘��)��u�A����ҡ�6v�^���`'g��.�C{q�2�qZ�{MJ_�LՁB4���f����/K�U_�=����% �e.�.����hԒ�Iy�J�xœ<L�l��K�m)1�O%�Ȟ�^-�s��Q?ie����r�e�⚐C��*�]z�43����r��w�/]c�n��:����Ѯ͵����%�"�����½�IG� u�y��/�2�>�U��{�+d��㢠��f�^#'-��.��"O��w՘
^�����~k�>�A(��W	sn��n �}�f�@�:�s�I�r��Q!a$���F�Yw���4�mU�ݘ�5�`?��7H��Ԃ��k����}�D�Hf�<�:��Ӧ�K��5/Qi	R��r!�(�Q�bpg���]*ĵ�WB�@��b��� ��,�k ��&$�7�����O�z�N:pK�Ei�C�|9�B��a�fwND��2�ҞQ�B���5.�e��T���c�����i��+��x�����f#^�%�+�wr�(O��!<������MQ#���P> �l�����!��h�2�N1Á���f��EF��L���66�7�H�{z�������f�|ɬ2/�W��ԇ�*54d63��%W��|�W��鲢��p�A��\n��`	����D�άD�o]Qkg�zj��j�e�ZF�6�Rdt������ M̕��p_Hbt ��@y5[�>�A��͵��~��鋤�'�=85^�gl�1f=e�L�h��������!������&�4��������`g���XV�ȪxH�g�-�(��K�A�⠁��5P�ʩ��9�3l~�����W;{Ť��h���';sj��p����M���ŏ�6���D�Th_�7ר05T!M�e1�ゲ�V�Q�kHxQ?�ٸ��g<���o��#N�R:��P�l�E{��"�+���i�)��m� P��3��<�{�&c�֩{QYg�K+���?Йs�)=z+٘��W�QD�o�ֹ(C��$�G���PZd@o�D����ʙH8d6�5Y��+����N���F����4�?�h�>��n��&��+uTCS�@����|��r�ೡ����j'��6y֑Xn5�G U�L�gr�|�\BI�,�$�'=<rt��U ���t�;�=�-x��9��Ntw�	U�zǖ=ٱ0����c3�e�f��h���1�9�^����1�|T*�lN:B^j�;W��.��s�>��(�<b�J�J���9�Gٌ�\��	��^�GU]Tzq٦���
L+?.���Cn�E���5;��_r��k%����L��bt���^*�����t0e�v�ek7C:9�a�wV�]��f�0���$��9��A�|��	+���"4�֥��z�c�̜uw��L��7���$vu~����;�03