XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���_0[kߔ�vٶfʼY��s$���n�_aUY��)'��������aGf��@�q_��dm8�G|�=s�U��F�6���Kߟ�C��%jaGD襯y"Ԭ%���
�t0�p��lyob���&�;-6��ki��9�7~m[��=n�|�)�
�%	���H�K��P�K�[�J����Q��p��2����*
���'MGsB���L�oV8RF��Y3�����Dm��0�4��DVe��MDК$P�<�2 �nh2G�犕���:1�.��㎧���`�&�eQ��N�*�mլљ��c��8CV�:���|s'+�J�|#�~BC8(��`��ۗ�Q�Ht���z�Y�6�"X�λ�����\���:�!�ʌ�r��$�nf��j���d�D�j��{��o��N��E��r�_���{'zRu�N��-��s$=�\>C(]�s�ȕ�{%ڴ�N��q��u-�i�])��o<��`P�m�0
Uc`����V�^Q�5�'7	�ZX�U⭌���P���M������p�P��9�`���r�oI�h{�����l�%����	�u �(�J��A�ך�ǘ��C_�G���"�0��T���3������P����>,�8�*1��l�2�|h2�*�g�tMuV#DG������k9����C��+��\��L�7�Ƴt�^�YNÙ|�z��v�,�X䲬b�2�����1.��eRa����A�YM�{��q��j����,GX�XlxVHYEB    39de    1170�2�]��_a·������L���\�~?�[.�q�^����&^�h�t	|�Pt�j��iJ�*�WO��ug���{�Vl�W�j�d�TBp�e��n
܋���pݽ��U����9��q����׊9��꘡?�-~1��7x<���r,^�}�Y�so��6���v3m�O��mI����!��F��u�K���M7�7YN>�3�.����o��o.�|U��`�b��������1�H����Y���@J,33���,t26r�/����"4�Ӽt\0���Ӣ#��6^rTw�$hf�e����-pd�����n|�d��<bD���M�_b��lg�6�s=ha96���$h�b4�q�����!P����^�	���bP���� �g�����3�i��]�l�2~@�u{S�&����b󡪰HĖj���?������L3b%�F�Tż ���d�AҌK;�ړ��
��2�y�o�x	q�-�`�W��F�W~����ȸǰ�U�J�R|��#z��@�5�/PDγX���e�@��w���й�M�?t�zxƀX`� ��>��U��Þ��'�썧Hwه	�,��ȏP1�^)-�^�@G��<���,��_*�4�xF6��2��Ǳ�>�*�w�*и��Z���y��g��QǴ��L�m�s������1�!V�hͅ�J������]�2��垛���� p�aB��n�N���r*U�����>��z�X�B�Ƕ���d�m�?5)���/�"�=�g�gIh1%!��i���c!��A�d�	��HL�p�,l�e�7�0�1��ze��P
��R�:�!��<�Œ�Ĳؽ3�g��bI«���=%�����
�1 #�7��@ǉ��c�;U�߹��a19�*�� �V$9����O��+���=��,N��eL�z�]�Ŷ�`ȡKE���pdf�
q�l�I,$��f�X&����.�Q�Mi#��Q3Y�K����\"��"xgKD�ȩrv0��X�����'Фr~�s��
�y�N�:q�1����ż������z����y�&� a�� E�L��<죤�Ț v��тd)�1�����t(����PZ��b��t/�|��G�>�7*3�Fm�Y��lG���ؠ��g��ڱ��.���,���,`>�E8�K�b�G $�Mi��}�[��`�<��M	���fٹ�_�I�(�\V�pH�Ό�z��K�e*� ��
�u��ׄW��k9�},`����,���6���5�X_	��z�I�
��4F�(G6tBg��2ם��hSω��d�~���6[�u���
闛 �9jazC�4�G��|-�V&��-<�4V��T�VQM���_MP��㚀���DH��;�|�R%C٦guG ��D��{;�73~O��E�"�0�D�b��}�����d���=��/�{���6v[�:~%�≌-�YkN.�	�d�@��0n^9��a۲z/�v0�a��BE��fE�0jU��y��``�%�wo��'M�ɣ��p��{Rٸ���/��*�`qW�.,��=�r�r���mQ
�%��+��g}=j���_ �ӯ��A�����������*��#G�2��B�1�.{e��O�"~�%3#T�n�=Ҍ������>�Wя�i�f�%q����D�6��@Ǽ�Q.���c���X�ߘt���cOyF;j欳.3 TvPߜ�����*�C�B�g��Q�޺\N�/<�,��X~�9	�����Y�?e�w��I}3�<��\��jk{��ا���	%T�s�`˸��@K'<�P��W����aXJ:��N��gtS�OǨ����� _�8��)�/���3�H'�Τ�5�,́��TIN�]z�5P ���o��T���h7=f��O��<�68*&L��ڃ�.U�0K��gz�#D
^�3��Y�a���$� F�Ǿ����^�ӏ����)�|D���Q Ќ7g�4E�ŻsM���_c���}�c�X�fo������3?K�M��+������t �Y��`~�j,��eq�!ox�ǈǴV�����OƇ�aV������j-B%��8}���hn9�����ILӳ�}�0Rv_�z�g(4r�K]$*E�M_�Ui�'}W]l>�74��~h���B���pCX��֧L�&� ��i`(�l�im�i����УR����7��LE�m\t��c&L�,�m�2��$C���{h�-cf���*��ov=���:��ʑz��>Y�P��m�a଻O3|�z��KC���3�߯�Mz�d���`��t�'�Ac7�ׇ�YsMW�V�N��W�SE׆~2�E�C�QO�|��bP*���HG
���+��Cj���C��4�\���Z�UM���$��D1��#�;<��P["�1.��*�=��%�z �������������[ni>C2�G mX��k�l�K7VN��Sb�z�-��c�`&CP��27q��EQyrgs�����0i�t�1���(�2�)/��$���/1≈�z6ʀ�O��RF�����Z��fm����H�/�GHX-@��ON����RK��O�Z��՝��j&L���|1���0a*Czv|��s��r�y�q��Q0���FK�?�얚�'��wb����%:�W�� N��D/�{?���)�EFN�D�S��A1�L�͕Ѡg�dW����D`�Yuݷ�}r�xu|�CWJv6s���'�$%�pBl�D�.&�Y�i��g�\lݓtP|x�|��>�'�ց�]?d���Hxm����A��f�8���@aơ�S�lu��ܣ�ߘ�O���̓_Ac��8�3�%��F���^:���S�P�Jo�8�wx*d����]"ڱU��j����~��%%��ߢ�a`Cu�f��#\�%��ҳ{q�cf�"e����Y���6�����I����y�d��VB,?O���S�����g�P�� �g��p��|��I}C(�"�m�j�<���
���N7��x15	�a�/Vly��P�@t�.��-W
,�O�$�`�������m��݀�:_���,�`�h��zx$��g�+���s�e�j*n�W�HM���p�tN@r���GCUp�B�d���8e��qr!���;L�F�:O�-^�Ka,濋sV5���?\w��$g,���a/��%��e�]�"���9��o �uL�˪����9ɏ2/px����ӱKB����~f���!	|^X^��]�IMC��p=Hfm�@�	��>��*�R��{?��k���[�Ͻ���U��Hs��0>��nR�p��$���T��5�B4pE\.!ݹ��$��Co�(����d-h$��s%�K�%0!?ρ��YI�?����Q+�����At�RAK�0�A����L�!�U��=>phn�Y�zL[8��5�É�H�ޤM����b��6���$kB�s0P�:���;�]o�˾ܣ�8��|�q���s��?�O��9��!e�O{o+M �1�m`�ҹ?�O9�^���|�J�Ĩ�ںrCdz�s��XѣB���($�B��>#'�����8>$����@<,���Y1�ӗ��uN���ȥk�[��6�p�o)`Z�jӀpor�gŦ!�R���yT��J���V+#����ǁvQ��(��w[�a�ì%G�ry�|�[lhu��c<����0G�F�+�'Y��9��-IpOk+��?�,��F~��@��o���������ϼ��<�f��g��-�nkM�'>�1U��+�<�����ǜz�l��	+��mBQ$W
�D$�to�
L@��X�X�٘���M���h�
�7�^%`ld�x��a<��<��+���b���_�]����P��$hT��r>n���ZW��@�	VS��	� �2i'��X�_��^t���Q�����r/�iM��`/S6�V��O�껱����g��0�˲�(9�6ʤ�Ř��a2�	��ޘ���#;��)���+9�c�m`xE��S��d�4�_�Ɣd+�ȗ1(���,����L�z��	���&]�o���dI�n�������ɤ���= ��1*�N��&
T�؇܈F!�u�LE钱)�m`�eg����]��>'?�S��Z0`V�b_"��f���د}��0������M�C��5Z�����9G�G�/n�T˪".j&˅����_��(���ӱ���3,����6��j���j
9V��jX�$�.�w��#���P��?C܂��R�H�]f,w��Ҥ� �	x��ε}�]k� mW�l]��p�c��୳S,�e=��CqcBn��9���i~Utݝ��@�㗕�	��)VzL�n�GK�	k%�Ŧ