XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��IV�b2�
v��e�$aW��.��qL�Gk�"8����w쇏,x< 7�2��T,��mI�a�u�n�:��6�H� {�VB�ﳓ������lP����c�&����e�|�)~d�'g�z�Q3��fi�@�3R�	�>�˧����ݩ��Q�ӂQe�M��F��x�Ĉ{���|���W�25���e�����n�L���("D$f;.��aLt%tfP���-���q���sYz�n�)���K@`�V˸Q8%ԖS9��_��3E��J�y�9{n���i�(�ϙ���1NK���4��0$�>3�`�bVt���pQcn�%C��^~}2��ra�׀�B@�r�.׭	6���_�Xu�g�7�����{�P-���PԀ7T�O��dKU L����Z����xF��m�;�"�oM6r7*/����+!=|�:���o]z���>e�ՋE��aw8�|^uI_�8�\��Ee4�gp��|�R=�ކ�e���[.�b��d�B�#�?�ܑ�blnJ�)����e��A�n�ɞ��~H�;�-��[G��|�U�)�#2౸���E�=s3�.�c�xw�^���pkN+_l����Դ��!?M7�nv�OD|��Ԉ�Y�̵
�X���d��wY�wf�yqvߏ��'r����z/v����6���B�dg�l���B�Mm%w�JЧ�#j��b��c8AL�f��y2��y�Sǂ��@ͱ��t���ٱNP=��3%�!wvF"�8Jd�IQ���0�|V�XlxVHYEB    28ae     b60d��I�E�S8�B���z�3ʟ���P������G\�l󪾅1����l��S����� f�������I��=»���K�f�Kי�B-i*}�y�"�>�(�1;]h ��c@�¬��������2�LF6����[(ڇ�d��ٖ@׋�Nҋ��~��r�D5�P���{�
�]Kɭ��Z&2��~�}�=��{�+��/����m޼er�䖵�!�?X��z�PIRH!��L4F�$��1"�g,�����5�'Lj�͈�&ȊD��3���x��[L`:�)��p��	0�u�|��,�D�Ϛ}s�U����:���a$pH� �������ﻴ�,���ck?����'&�� պ{;1���*�j����-~��\k��9��&��@�N(ǆ������W�����塩O�YJXKd\��]%Ĝ\e�?��7ّ��d��c?�#'?��%8��-f�{�[�8�]����w/���@">E���C�9R"�#I����)#׊j�Q+vA�jg�||iyB
=�jo1V�����Pm��q����B:H��)(�~n%�	�a��v����������]�L�eˀә�r/�k\�W�ߎ9����l ����~@+�6��Y=�/+fZ���=@�v��,�JG��N_�/䔊>�A�M���ttL(@3�ϓ�o� V�k���-
9�����\� �&/+..��7�*:;z�O����bNe�"Fߎ3{t�]ԍMV����^��oN���Ţrhj<����kw˒o��*�����vp] )�$��c�ϸH�����-���v �_��\��D:�ሔ��NP��r�D^�	
z)A�A0r��8�11��[� Z�A$EǪ��n�;��V���U��u�{����~к���L["��[y�Q���%x�|N��B/i���蘺v?s�A�HA
tF*�
�K>_��QR�3\%��������.�R��+�� ��
	�W�j��߾�f0'�ڳ��q~7.�����ߠ���x�����)+p�6�$�С;3���v��y>Q�iRg�I"��z��(��e�4���?r�C�B�}�O�k�s�*Rڤ����z�i�-9�lovY�~pf�y��ّĆ��֙�"z�m+�p�N%.ղh���5D�U�y���͖���"J�0�;���w�Ը��[�õ�������r�������,H��"�I�s0���6�g�m��X���}I�0������n5������y�G$����^(�T`��l1��a0@�r7;�b.��%�Y��KK�8؛���Fql�xMnq�Bʡ)�7ٓNu9�h��]�}<�
/P<+�ݣ��s[�ű<�Ǚ��y
k-��W0����Տ<*~�hن���*����.�\�dgx ����LR�\/J[JP��X5H�(7�:K�=cs��	j��Y1�`h�o�e�S�^d�2��o,��%�i��z�����q��#��U��웖�v�+��%	R�nU�'�f��Н'�}��/q�h���\'Y�/:!�s��&�Vl���A��<�_%U�F�!� �j�~�����0<5)�8j쥉��so��^b/L��ǤA��n��i������$w4�Q���O��1�DsZL<0�<h���n��ģX	B�P�l����-%�g:�	8=�J���-�t	�6�^���˽8�"�b��V��IȦe+<����H�H���@#U��{M�Z�9�"L��\2�
�&x���
Z~���{��� -��7�k������dD��� ���V�����@] x>'��)>��!^D�^���gt���PD�˘O�!�$r̎��')p��y����\�?}�<��S"G���J�����0Q�%��_^\�ߝ��� 
�	�χ�sE���5y%����fᑃ�E2���6����}qɍ\,,�e%�w�mo��τvBTF%Lvg�I2ҁl9�漩"n�}���,[����;�!���cE�Q�3�$�N��p�F�8���y �p M���[�N���a�H��Z�D���H�Nu)	{��M�*)l&S���_|0� [E�4��R��$���� �Y��� �;8J�c�ex%��+q�gN��1f�XFx����ˀ����?E�cm����'�7=���~�ϔe�� dP��Ӯl�<�}���;\z�w��Sj�e(�p����P)��h�Jn�8���x_-̙!]`�ũ�gLz�Dp%�y�yݑ�X���,�t�7@"�7}i�Y�=V������&�VE Y)�W���jtL����|Jv)��O~%��M���7�9��i[�K+.��TWE��8�Go�C<�H�Q�>�<�X;�5g��f�A�؈U`\�����k&wl�F��.W�p����⥉(�$΀	�6NƤ��aLX��F)��@�UM�$���SGQ%IF�םA3��GE��ا�˥V-�L�v'������##����=��/�����@H���ƐMr�@�=K�S<�`EP�Ӗ
Zl�"����~U\�9�Yb�/��%��Ў6xHyA�E	�:a����[�O��$��	��M-��:�׾=I#�h��|�O�R���Rj��h��_�
��ӫ���c���!�7�NV�SW��x�^u�ٱ��/Ӏ�Bu�g�}0����d�ԗ��M
%�_��dIndC��Z�>*V����x9�n���h�w^?�K?���8���O5(,�_:�\?��@F_��q�,qsI�C	�7v�y�#�b�	�X�t� �=M�F&-���v�j��Z��G��voh}��Qc� �j�+{��	a� ��0��7���_��z������:X�j"���d��I�@-�Mx#��v���|�.���W����1z�.��