XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��\UU�/kI��>�ږ�Π������X������@sIs����"[ہ9x�GE�m���iM�7�F�z�> #��0�!��s�����!X9A:������oz&�x���(t�e�k��6Æ�4F��o���&|a��v�5&��˿H;���3���8�Ơ�J'Wʔ�圇eq+�V-�@[��).pS$��!��~�U�֖���Z��`)��n�3[iV��ྲ�y�(��e����������Z�>��S5�;38�2L�ܧM\8o�nk�ܿ�-��yD�v�$�o������"�]v~v��O�:P�U��+�za�a!]��G���E��q���J�O�����)	�-cc�����|W��mh[���ގd	���ߥ�jm���6�l�u�bW	�f��OI��wu�=���BZ�2�~\B~���<� �%��N�ª�.T��D�Ԅ��S�
��p2A6M
?�
�����nX/ �q9tY+b^���7��8y��\62y����ޣ����W&fQ��&���ni���>eD����7�n݋<E�$�E �$�I�Eq=���4��`R/�L��tZ�A�\��F�)̳,o�H�s�'��&�q�y��L�1��_5����Fln>��/��+����Η���`��L��_J�� ����p���7�&��򱹴��In�NGWOXb�{���Gw�7���	��i��"\ք.<a0���i2���K����B�ء-�K-��f�0XlxVHYEB     e07     680O\�|��lI�~�<���&�ҌP�����rTч�6`18V?)��I~�H��g���_q_�Z�qLy?֧*s���{So@��ݠ�N[y7W�����5 (g*�]��K �T�%S��dȬ�����u�
��c4ߙ �x;1#�-@�|�	B��c���p�F/J>��`0�Im�jg#����*k���:.�}h�ao܇L���!����vf/�/�����9j�4�XtW���[�iKF��Q�,�x�:6����Ot�QTȮq|�"q ���#r��r3��Ix���aEv�GY��N=�4.�	��j�.q�B�|a�|+��k}וq�d��/��x�`_U�>�7����!��:ņ*������e �[�>¯����!�9� untb}����=�"��a� k|���H�]�b�H�¸�Dw�o��;�Qh�yK	��%f{���=���m2�o<��P����Z���|�Ww���t��Ӏsq�� �Z��F�uK~�1o�,������j�r%ǿ2����5��m���PR5���Q�+gnP��m�/K��wӸ<8-�]�줻���O�i�Dq��S0��V<�0��.���ڂ�ht��P�Y̙��*v�2�=p(�Y�!ݚ�D�uVh�<7��<S f�f��aƦ�A��W%����-�P�*��BБ�lT�����/@������/�����1�;�Ncr|�
�}�T���v,�L#�}>���~���kK<ʄ>QA�d�@wG�/6�n��o�2c��盤1� ��x93��Η�Wr�~�Y�~�eA�?���_��Q�8ɏ�R$�dA�!��	�����l�?Jk���b'���s�m�R%A�+C�4R^��C���/M�},�ߵ��|����A�}7�s��������Gg�� ��Ŧ㫜H����(��_�dw�#+9�5��MO%�`�	O_0i �D� i�]yx����b�-��ҿ��.��[�}�̿�ۤ�୪s��!f	�q虓*\B��fwd�����\	-�.Y�h�k��C�˱�b�"��2���[Ӎ��wh��t�:�-<&+�$��4S.$�&J��tH��`�1:�&MI,�Y��*��¨�HVeF>h;���JQ�����Y ��[P	�q5
n��,2�:��Y�W������r�hq)+dL5_W����S}¹���|Z���v��+�/��՜d���=�p�
��ɠ�)�׈-eސ�R������q��-���O��u�o5旉���Q!sC�mW0fv�5�w߀�)�g�y.�3��U������:x�S4Sc� ��zYu��i�S����d�+�[-�Ƶ�&��Q��*%����K�  TA֊9��\C�|��w���S����ڈ%-E㙕��O�B`�F�x�\ACy�y2���� *2��/ø�5����rS?n�3 E;�b�qyA�ʡ�'!�����M6�3b�7��9AK��i�q6�6�S>���5��Ŀ�{�'ߨ������$D<��@��f�"�=VT���X�p�1osKsQ����DfZ�{FTH/q����
�O�fA�l=�A��m<Thc/���:��� IEm�ʴld��ⱛ1Y��C;��bρ+����u��7��CX�P�v