XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� �W`�t�U��z 1	��u�M6�,� ���
ۑt9w��^��9�KGl�����xg��X���&A�6�=�����w@~]��$��~H�q���̃� �0A_CEő�n�䱈�6��x\���L�t'p9��p���-Y���[A�&O�&�7��Zz�Ѝ	�՛���(:��l��~	K
5�N��MX���SFW���ϲ��1��v  Sm�jt���Xij]�ɗ�B��ي!�l+08f�3����b���B����4�W`��[�P�|��cz�R���B{z=�o���k��=�F��NO�yl&~]{�Z�CZu�Js  �X<O�>�p4N͈��{��n���~�t{;h�峂��Z9:Ȭ��Vp�Hz�77��c��P��͉�?�l�C�\J=t	�cj��+k:��J4�S?����'�}vg�S��>�Qn3 <�I������+gy �xX1�<��%>�o�"l��Mb����zҊ���ᩇ�����b�F�Q��nꓙ�K9�}�6�a�Guϊa�>�n�Y:pgÐ"۵��?!')2�
���-��W�Pk�d:�_�G. �G=��ɕ���`�C!S��ꋴgV�(R�cx�u9م��WIʃ�O��)��D�'2b^�IV�?C,�l� eJ�Ń���\���{�'�*7X��ap��������e��RqB$�2�t�<׵���d&�+Z��o��@��� ��y��B���n��- gq|�!�3ծ]�m'���g�
�+XlxVHYEB    1ea4     920P)��(O ���������KĘ�Ȑ9.�;������"V�Q�R,�7�~ݛ �_�?�zbUm�7:�D����J�XOf�щ��]�Բ�o[s�p'���qE���-�m���зG�2�vdز�p� /�؈*�$F���I�nL �N�cϛa�������β6n���Y�0��K,k��n�OP�@�����2����T1�&;xA��W��O/ŏ�kV-���"~�Y9i�x���vG �N�C�?��-�aO�C�L�V9޷�|�OI�i�:�(���h_�ؤ��ѬG+�"a@أ�sUv�,'����3�4	^�9æ���w�#,�7-G���h��=_j.���
Ǩl��%
�5�=&��������]�~�L +-�_B ���#	h}�v=V)g�u�(�о��|��<��^e����߂Y��Ԭ�8cgNio#�Պxr/��93�Q�&�s�������
����$G��/f�����׫�>�s�#�_��k�P	�\�A�|L�u���Y-̣��0S��}�V�2ry�\v��K�В=fkf�O��S�+���r�i����Wo�|�˕V�4/[�&�DKQ�	5_)�ͱ���ת=�����r,�jD�[J��U�j�g�;�A@�yB���EA>��)(<�~����l�;�xG�XJ����M�jW� �@�ˉ�.,T��:��j�N.V�A<԰�T�#�,�%a����Ͱ�&�?C�J����O=���4�K=�e����E�u7�3\^���r�@Jf�Bk�1��!۱��U�Ӄ���~���.IU{�',�&E�l�~��٤f������>H�q�f�_w�бׯ<�g/���0��OS�u�ƛc����5I0���un���i��5�9��u9c_�����H�M޹���{|;��C���� p���p��0=״o����K����eiƩ�|�lMY�d�r�\kh��Sy��(��N��l-T	�
�&���J����z3��u|�������Ejd��ϲ�6���LcfQ2=RK{��a�_"��	�$c��Fc�9�����V��I��0��X4"�I���V���G� ��v��<��G�79�b?��Bɢh�r�z���:R1#�# F��&�{� ���e!��o�K���� �g�2g\g����)���
o~&{�8-��L���HO;@�.F�n)���o!�������;���>��BVF�9�)Ao6�\A#�����	=j��W�ac0��� ���տ�^0P�_�����C�/Z�8wi��nN+��7���P<���n+k]����"J���j�nn �.z�zO��?�=~ר�R=�� �_ z���>��w0kNծX㔗��^æ��7������h�E�%U ��c5���[F���f%&Z����mi��1EO��f^��qnMQ����B%-�"��=����!!�s��\ϱ�*�ޤLS˵fxT7Z�Na����I�a�bP1.gX��o�7�q��[��"��?����\�y�	4�*��8Q[|�`�rM�g��N83¼�k��^�2�}�5��VfS�+�i�����YF�0z���-&��!�/#N�n�(E_�,�(��H�RE7�
��zM�n�n�-�t&��ɷO|�.MW0�����v=*ib�Z�@q�7�����j��S�Kܱ5(yC�P.��X�������4�r�q����b[�%�t�k�4���d���!҅�Z ]l<��S��8G�n#b�r�#=�>
���̷��U�Q��=�t�`���;�q��B��Ev�!��3GLnI7E_��`���N�g�@���D[��j5�ұo�L���(%^�}�=p��ط�A��U\{��؆����~�L���l��|ק7�;��8��S{��f�j���1���/B'�-�=a�/03�M3��@�!s��!����fZ�U�t���w����_�M*l76��ה�u����L�j��uj�f��2�Yk]��2����j�S�dڈ:gX�H�H߶Y�G$j�NUT��۹�ޔP3Ox	"����v��ɚMUl&ZH�U�PI_�>��\����#�����%��y��/,{U��]�������(~,n<�ӽDρHb�j����ui	��;SdP���u����0+�"���/�c��4#2�4k���p�魖��\�"�&#,�����_�#���j��2���ܪ��Ȳ��e@B���~؜]S�t��6��'᛾�`�L$L�TN�L|��T=CX�w�/ő