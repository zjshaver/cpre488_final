XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#%������9cc�k��7��/�GԂL������vn�=���c0�b4��`�{u�	�V�l�C`����b G|P	�ɏ����R�����	����#�F�C��y�=���jMh�-8�!�����������؝�>ֺ@����.�˂?�`~���d{[F��XȤ�:	4����H�L�o��&���kz���cgHqp���r�ht�h1K��A����ߊ�z�Ǽ�S��ց�|�����\sr����ښ�,K��|c#�
��brk@&�x"��]�y&ބ^��U���/b�|o$���TrQ�g�Ď�>_��n����h��N���f�0�f3N�`���h��;�q�`BDw����
M���/�&���ݒn�#�������Ͻ;@�,� �K�.r����6�9�
��.����X�I��������^��m�*Eq���֫P1G�C���%sO��]�[�"U\[SU ��J���{��N�'�f�8"��%u�����a"��I�et��M����2S.����֮d|P����e�#�#;����!C%��2�E9�����`���وBj8��o��d�\i.��6�]t=���jd�f���B%U$J-G��}�	ɄY�=n��m��v�-���'�-�1u�H�B�� W~z~r�oV����/�1~�v�8�.(+�1��{I��I,X��I>-����¢�s���1#>���y�C����ċS�����d=���m_� XlxVHYEB    48e3     e00W��-}�9�m���Ϯ�	A�f��/�v��,UƏ��\��K��(O��9��O�����	�G�R����)r��	 �iG�j��pX;��a}�ܾT�ΐwب�잷Ջ��(��]cݜ[x�Pq}�=��fxR>h�q;嚓�=�� 
�lM�kv�c��\� ��S�V9|CA�YB���)��`��rPe�>`q�S����dAG��3�� g�
2f���u'�W��q8���s��m�;��ݦ-�#X�Q��DpM�|��JL�����jc��L���7��
+dV��$���.�?��Ķ�o|�6f��~@���n��D��a�_W������1�8�.�b�б����%��5Dxl�\����;�������) �'����@�q�̷���`���v��thm���Wn���F����ԘR�mk��6u]��#nx��"���) ��H��:�Ԇ���������4|��y�s��i���L��u|E�b�1h=��Okß�vo)��Q O ���4��h#�N�p��qې=(TS,�Б�Hm_]�e�~�+���h��p�V	��vG$"1,
�>.N��m�����q>T.%��6@J�k��JTS�`�L5q�Rϙ��6\���Q�#n���*�0J��FO�:��-�ŗ`�:��a��+nK�U�=�;gO�����������KvE0r>���t1?�с�@�z�,%�us������1��K!,��|Z�&���W�v�J!A�5	$d�g��L��B2�@�H�!bӀ�`�*fM��_�-�¿Ɛ'�q���[�R��F��8�_Wp�v̚$�H
��°}�dR���|�y!b#P��`�E��;�!�#GP5�&$S����������r�!��{��	�"���\֟�$-�c�sz��"��*��h('�]i|҇dܗ�:�ʫ]����f\�
�����3�IŎ�}�7#�¸α�N���rܶfs��t/����b��#4�AƆ�&����x˵m�#+pWc/S%�J:����òϬ%UJ�����s��4tGߪ�>}�ȸjW7�v��PO+�����D<ObE70E
ժ��\� �����J�w6n�oE���O��Q����o�������@j���C��$��Q�m:�����՟�7��GF�5������o�S�5ڝ��W4���1�G���W��L��y�4%#c�޷u�,��^�kn����4%�5ML��BG
�şյW|��ޭ�R��ѓ���hd*��������(��^�f{8&�vP7�s�G&��Us�~E�փ�k�%�U8������m�����:u�r�J��o8����MrG�v�Z|ge�ڠ���/�mV�`my�Ьw�1�g�j*\��J����|�&��%pAe�ZK��!����4��?�,��8��.����z�$_����@jxU�yr��&S*��p~5r'�ʛ��G��w��������M��3ul귵��1)�0#I^QkJ�c��ϵ,a��y�� �3l��w��@�̨5��+6������U� .��M!��Yv���1�G_��!jN��B[9M|ٜ8^p�۟���<W����=�c:�,٨���֟�:ȡ��ȋ��	��Q����-D=E:|�GV�#+�[�T��`�@:�A:c��Fl/O�nW��5�Z�E�x�2;ޥx�l��%4z{��WQ�_Rz�tT�$#���(h�,��<fê8E�!�RrxT�\hߴ:��PM��"�ܤSOi��و�c%���K�ƪQ�AĻT���k�s�uG�M��Iu�V�3��q������et[�}����{L2�������z	������ɠ�y�:�����$&��c�Ӱ�n�P��89�����h��D���*�'��+�EL教�Z#8�`�ac�����`&h�3�娞���#��SJ��-���#���C�wn�����"��k'�0���bϏ�M�9�^;��*���裦E�t�[�(7[�y��s�΂U��F��*q }zJ�A�P�
��Ht��@���3�#��c@B_�d��v��y�6�iJ�>q
�u�m����:&O��[T�fRɠr(�w�ee%�(-lƝ�'��!��3���%d=w��Y�ٺ=t*,�����4�ŭe�e�7��.!p�觪�\'�����Z}٧YUv�4�I�M|Rm�p?�]��
�FRXH�aV��42������yPY�2�.�J_�-Ow>A�g>[��!+����O�n�����avA"�Ϙ��)�ZS��&]�+q@���y�`mov��\ႸZF�<��Q�	�F=l	�|$�҆D���j��ȷ�myz�ϗ��հ 8��܊��zrnN�U�t[>D��������B��V;j �Km�z�G`���=�r�I�?���QK=�g��Xޟ���ͱIZ�hl�Ns�X��c�ßg��S�tdGc��`L���Y'UY�����V8��7�9��kN�-��X�vu(q
ZR9i`Z~��[ ~R�G��V���s��\�\{���� *����`^����/l�FWn�2���ڝ��D�ܲF�.����c�/�{����Ž[�`���کTY���nc�Q)W��؆��*�%I�'ߪ9�޾�51��^���!���}ĊĄV9��1��X�әn'����H!��[0�#s�ux��:�n��K �_�ScB^�+I{���Ƕ��:NSZ�g+�#�d�=� �+:p5�확�����ϫB��E�ez�t�dB�v'zҩ�Y>����u?ޝ|ᎱU<�	DKW�"Y��C�(� g�[�뵘咾ma��xa\R��ܡ�Qv���s�b��#��d�$iϯ�噇�F���=� �DE�����7��&�����v�*ݤ�+�͈O�'���n�� 氅!7��Bґ���T@�s�j����9y��F.�u�}��vP������,����x��8U8�iju�����������Ơ{	A�$��)8%��TyKa��B�QWe�xfb���Et�}a֗������3qY:�Ԯ5��X����4[Qw=F����͍��X:d�Vb�/�7��Ǘ)@���g��ʒ�3��J6�8n'a�����d��]���W�r�F��'	\5�2(:w�wXt���f�.��n}�h�S_[����L�IV)U��심�&n���A���p����+Y!�۩t��gʿO������E���d.X���S� *8)��Y��-��	,脋бW1+�K
��|�56�I�G
]�n�f�����s�_$���d�/�Jzj���ʉ�$y�^UI�4w���S38ɭa0*��FS��½�j�i��kc�@�Q��M���Y���.hZ��u��.�������ڒe��"(� l��x�F���-�,�pbo�)fr6Vq��� ��W̿v�i*�bsm���'��CC��O���|$�I�o��M(-c�rg.B�M:���?kf�����Y��I'����կ;D�<&�2-�����