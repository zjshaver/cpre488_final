XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��^<�]�UR5�M��}/��$��I�׆�����ȭ� �t��lfF5�+,g>�بв_Q�z-+Y�����X`��,5uu�����|e�}v#o$A	K��P���*�یP�����2k�%X�\����g�"��6���_��5�P� <��;���� 0��(�������fMO�('�2f)��|2��^�ax�˿ph ���{���?��*�bS����4�Pe�	<�CV��EgY�^�3�h5��,v����*w?S�ڞP�%��U��!�*wou�
Vl��S����hU�c|g��:��I�fb�	T�<4+�����w��g~��R0��!��\�%�ڥ��q*&&ł�I�q�	�"(u��pz��X?�:މ�cՌN�1`ޱt#�4�S�yCvSq�iG�m5WCw���@G��!�њ���F$��h�^��tn5�=�b8���еY8c���I	�*�v�N��x��1.��@jܒ�R
�j)�w�����Tݥ�ex�	��@�q���PS�.�7\e��!������f�>�Ɨ+4���(�����f5���W���^��9P��� 1�����
푕�a����M���0��'dc��K��&��˙t�$��>e|a ��:;��	0<(sR�9��	���T ��B�yŧ�>1b:=9�>)�a�����TR0��?��B�E�cj�����H���5�z��8�S-�T�K1�iS�h�����~vP��Gc�e�XlxVHYEB    241a     ad0W}����j9-��%�w�J:Q����EՊm�|W��E��W8���-.�5�\x���ǩP�<���*�@�(��B���T1�YGja;�ZZ}Z�0��Xݸqo�}�.g���Pw��GS��n�����P$�옲7�52�oM����~�8\2�qU�PM��ߛ������Q2<⅐����A��}��[��<!��
poyA�ս`�U������]�/؅E�C�n���P�p����2��C~��_r5 �&FpGU��!�\��A�[�Ml�	�]�ڴפ�����E!����1Qd)2�:���t6&��MD`l���bk�ú?v\�$���EY�� �;��4Dk��uFg_.�]���cC��pQ�e���Y�-w�h�
D�4DL�Y����e
��J��dT��_���	_��:���?�ˇ�A�2AC?D�rv�B^Q!�� �> |M�C�q#]������<������o������,(��X2�&��J٦�D������?�T��v�!	�-%.AB"rA�˨��`ī��lɜ96Vcے0Y3��;`w"��4+iUع
��ez��x��k�%�AsA4�5���v�e��dr���luRp�)ksI�Y|���C��o��kր-���L�)Nd�r�l̡��HX>Q�1�\S_]��0�st��m��F-1M������mZ��%��b���>�ƀ&D�	�e��� h�Tep'p����79ԔII�#|�
��h�V<��!Hu5���O��\��E�ʌ�0�z����H>CQ�?�`�}T���b���$�6�/���y�Om2>��5���wq�|�L��NP&1^:����5y�����B���YඵQ���y�x���i�sH@���S�^T_ٟ��@��ê�h�}GsP�t�H�Y�ydL�J5:qS��
��٧@�j���y7%'��+��%t�F�LY����w����;'Q���C��"�z�$���/k6#����z����|ǽ=�	���P�z�-�.��Bk]�
�n�i�9�y�!,2�'g�F�*a*#R����zt�}�4x��e/O���
&H������87��f��Mc�dx�S��!#Y�Ȥ�6�ҝTD��X�Px���������vĳ/1�qq�E*����W9�/�i�
���9ˇ�k �{N!x�4��Q��4� �����i)5R�����==n#i$2TB�����.J����t_1�c�W�&n��9�q�颃9��6$,9��_?��I�7�+�i���]���3���Np��%�"�bW�5�W�Sw���'�"i��-��o�"]�2�F�#��Z�4e�����L@BM����&
L�Sء��t�\Ƿ|%ʖY��7�	`�sz]��� a %n��Ǜ$T�$>K���0W���as��!�H����ͥ��Vc�[���XۆT��"�[O��ޣ�$��<�ש���aQ�Ie)� �Y�)pk�W���!@#���qh/��j��5M�>�[C@�ȅt`r �L78�F�&����4���>1j�JDL�D���QCus�e�`���'����P�w�/��i�J�z�{à��'7�R�K7��|�b�[�k�QS�%��@��;�7oZ6�h�14���υ���n�'���)yΜ���+�򻻺5}R6����הV9���;���5���ԕX�) ��;-�������$\��C�aR��2~���k�λ��+�T-Ds�m%@�(�*�k��/��W~�(�KR]��E��NX&��iPs�� ����E&?�V۲U��h�}=������痠��y~MGJ��R�v{�i�Y��M-UV)|I�˹z�'��!\��t���?e+9j���qkg!)oϼA���R�c�gkX���2�������L�j��eE4q����R���d8���s%�L
!ĭ/#��䂰-�Ɠm6��5+����$�J��ڵ����4q����� vYJ��G�M��%%�I�����`0�4��v�w�H�U1l�$!��գ�g��dA"G@����`Һ�0m�^P1��9��\m=�v0���k/B"M�N��R�Hn��[���h=ƽ�����EY�z��vחҲ-��f�U��!�X�'^�龨"ۢA�hQ�rJ�\sV���a�=ZP�L���%>��)3�(�i���a�*��3s���
�.�5�7b:�R�F��C^�:�c��a%K��*j�/��G���R���|��p e�r�E����21�t^\n���\P1�?��]�N0���[�=L���C����i�
��P��������k�6�H�
밄���0p8�H��BMQ"�×9���L7�.y�t�vH��k4]<��Z���
�i����2O䦒�ځ>7�$G���41+OH��_�|�T�m����׊A��p.��^!�a����?�w�#��,Y�^��Y`�4�����m��_�7�l�dh���@�-͗2|Ỷs�N5�""�����"��L{�"�9A�:o~R�J�M�Q^�=�lk�|�mۣ�}H��Ҧ˷�튚��*R�F�9�"�Z���d2����mǝ��,��}�R�:⮹���p�
�։�z��ȓ���_� t�`!{+� �c@Lc�j�(ɹ.V6��3"�N~��\x��AT��I�Mk+�;����j