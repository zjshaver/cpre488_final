XlxV64EB    5fe9    1830
V�4��W��%E�-~��}0����w.Pө��ZI���Q��I��czcĭɎ�L�:|�r�l5�~\�^=*X�K�:�����>��{B�_Dc�Ǘ�L�h�w�s6~0�ƿ�u��.NI�Kc�ڇB{�ε��xm+�f�����c��ʤM�w�Х��ݐq�TK*��s[�^8c���ýG��c\mQ�R���@�#�L��W�w�ҝ�Tk�\Rh8l��(�1�$�����_m�u��G�}���� #�Od%���k�.A�q�OR-��
ܾ��?��<���pX÷����2Q�3��V#�i�E��[��<E�b��$�5����<�)�x�^�-=?�s�ҝDT��j��D5�w���~� �5������*E*��~V�[��a͐��J��!"Џ�x��"�X]Z7��1~x�H��Qr^4�my@�*9�ճ���?}+��~Ʌ����8�)��^�d�lMق�sm��e8��F��M�(7~6@Oz�� ճ���eaP��M����p�j�OE2�O*���8�E�v�,�	�gH��rJ�D`�p	#1J�O��Ų7ӹ4�v�o��Sv9E�]Y<^�Ĥ�"����x��$�(z����WF�6�
=�侸�x �par�lٕlR#zU1�����\�����S����S�'-��ɀbgR��0�>Y9H�F߰�����s�����ہ5�hղÁx:v��A���R\������	� �^w�	\������~P�;��ǉ��i%��(%�C�����'�ދ��b��n�2G}M���%	����
�k�Yt;��^%����yU��?�k���\cic��-G��3��:ŧP������)W%�)"���Ѭ]6O�(��U?�,�G�D&�</sH�f�-�1 '���{9��Aa_:S�[,A2X h:��\��k>mp}z�K�K��&4=*=]%_p��
#ZdYYjW~�؋�Cc���I&�����b��n�~����gqL�������������){��3)��d2��ej{m5�/;�N��+�S��t$��G�SVy�.��S^�d0�B|�qfS�tWhrN���s�S�^�|2\v�y��8"Z��&Fc����t�)e�^.7H�a2,	.H�S��~o��gQd���x��
y5|5D�+x���Z�@lm�##��x��Ҁ�$�%:�~�
#PeF�bt�p�s߱��G��9g����"��3o#&%�sP��#^��*�U�#�˸/�kpL�s�_��]%��Q�;=�$���Vm�ؠ��/�w�/�F��&A\��-9��\�R���ҧy"�1 z�-��7΢Do�����=jn��p��EѴ�	n3l�
~^׽}9[+���2蠘{<���+o����T-���kQ��~ǅ���>���{��n:��%���a	SW�Ce�Dp&�[8�Qj]�~��AI���5�1g&�Љz����m
�^]F:���S{$�,Ek�؆Kē.K�]��O��t���+��1u�.��;�Δӳ�,�p�8�#���a0+���}�&�&OQT�ȉY��I4	!�o/��%b�Q%o�)w�[�Q�
߸�����=t?�)�u���C����_K�}����aà�#Ze�U��hX���4j25���y����T��KhR���h�c~�~܍}��c.O�i	�5�v���,��,�*���<�dBO�����`Ft��z�wȚ�SM�;W��,z���q�e��Mf'�7.➰��8�ĭp��6W����¯&5��co�� ͦ�z���O06dᘙ���-�g�x�j��k��4���^�D�ظ�ak���U����4+� ��[�-埽�q�$Ƨ��B����]xT���K�9��������\'5�JI�51n����"q*t�Ӂk�R3�����)X����Q!���B�-�t#m��q*K;/�֟>��|֩�=�����E,�>�]J	l(�0���kSĈ�pR�Q8+F�� ��-j��k�]�᠉�
gO�@~ַ ퟇I�������O]p�_������n����42�A8KmD�@��B>�wW<�m����O]�dYlK\�A���*���d''^]9���<��j���E�lƋa�m�t�\�?@�K�Mg]i��Z�-	ͪo@7�I�
��c�c��}=!�:�SR��MkK���W�,H�<k�d�%$��e����aoē���z������O�N	�D�UB��8>*X;U@骱�����>[��ðGƌJ�RF���l�#~%5���@�2a {L����l(�?Zø����Z^����� }��p��I0��ІN-��b�H��#��d�:6)�� .Gn��xw�HY�w�ȣ(4��>\�?��5HĘc�rŽ�2�ֵ���g�PA�E���W�~$� �1i�)���E{;����=�P�T��cW�f�:?�.�@Ք"e��	5f�q5]vԆM��i2���z^�!�I! <y���JX��6�2��}�����X�\Ǡ�6���!-�>v���h�b�wM�y�E��Mx
�Hjk��vl� {V��6�b����'\ŗ-��?;J���L�����X��x|���h�}'Q���&�Ѣ�ؿv�#~GA�t��B;�>�5�v� 8���5���E���Z�	�aa�t(�����_`Ϙ<��JOq��C����D�t�=r�F�
$B&���w�%�o3 I�.ɪ�d)m?I�R����B�ǌ����ao'�CҎbWOAHέ�'9E3t��_Nd���eCZ��1�вXl����`ʡ�����K�m:�ߜ���<�ȷ�d��2���>�>c�E�~19��R$fP��j����L�j܂�[T�j�?����	\PǱ�t*:����[�M��7�i�������!
w>�7��Q%՚�����ӹw��Li�12��<`��F/7�y,��%M�YG�l�)%�VϓC��tz�r!��|?]v᠗X�0(�����~ۤ�j�>�]E���%��7������+�q��gZ9^)�Hp�ɘ4�$�8 %2��������_+,��p}���������)�c�b�Fo�ɟ���c��ڴ)	��=e~������K�����_�9�~��ޠ�ǁ���&p� �%�1rdX<,wG��5G������sډ'��ߝB*8���K�M��"��N[[�j����씉�ҧ�-����3q�͡p�q�L����������2�=	a���5� �膚3"���2`9)��Dq����y��3�z�3n$�Qvڒ���u���d;�`R)�"� �Ԙ �2�4�k�|����h��k0Sش><疛F>M�M�����Y�S�~׿�m9���T��k���8>�.Z�}�I���CN9��5H�1h��7�0�Z�I4�0|�Y�5�pu���� �UH���#���P�@��Ó�.�F��֖�%W^�Q���sU��<������
V��P�lMC���A�c��**)bd4�8�S>6�V:�E ��&�:*?������^ c�1ɫ��r�?�� �Êr��񓷔Z.�N��@�e���^��<�'K�Qގ���ZG�(�4,W�a[ԋ9�rkk��f���'�F�
����Ɠ��U#W���"0s�*D%��/�X  	�x�ȱNy77G�c���z��7�S����M���~Ql��\i�9�f���B/���j���3Ռ`��-�2����^a�4�y\,r_�Pb'�)��I��n��;�ZKn~kР�es^��1.�C��J����Ҷj�⹗��UƱ���@��x�;���椵�� �zzZx�>O�ƈލ�/9)?n-���X�;䠊�N���1v.�q��/�Ed��Zyz*��E |��譒��(EQp�����.���:��/;�+��Z�D�g>6�=єTf��<��1�24��a�0�:�i�ͧe/�&��q�
^:��½�~�ƴ~u�[�x/F�n6�xc�?�����1����%�e�����	*�ڂ�L����~9l�؎e�%v�Ӳ����YCI�c�d4��:n!�j_GH,�id�)�d���qg�2�C ��҄�>&����	֑^��Gqv#w^y�䕌��U�!T��h}����&0mӟ�,�d��w�Ռ��9]�!4h�O�U��K���.��H�h6����;˷����A��:6��F}���QY��Pj��jv��&�@�	�p�x��<�o��=�|[�o����>�]2��3��Vb�[��q�)i����YF\��"&A��d %sξ$e�^4�;�tĿE��Ve��Pif"¼͝m_FQj�4�W`}��2c;|��7?}�aϟ���e�TPZ�ӥ.��j�(�����D)r�jG�lm�Fu���]cM���4(_��o�_ͣՍM�d$Zbq����Ṹ�]��gV�S%�d~�~2F5�&<��:H?���`ro�Y��i�}O�+��E�;y�E�͞���4f�����K���xJ#�zn�*�*��OX��lf�;�o]��E��#p���"�g

6������Crm_�(Q���iGٻ������
��\2r�?����!�������%�$����iz�����Jް�)O<��Tg�ln6�Z؞���$0/x��禊Q��ŗ���2 W7*�'z������0��;��_�ĩ5*��C�)�qG=_)0"�,�)k��\��J�r]\�89�}֟�m��R�劤��%;k��O�5H��@|Y���ѳ q�ᰰ*n�/{�Kł��vB<��x����#ɭ^LO����ݶ���e�de.�`pF^�`�����uB��"~f��<�%�\1bc'�Dsk�[�fWJ���0:]�`TJ(��3���{�{��$�q�{��%�lOڰoļ����\o�p��G�w��;�<1��NY
�����⪸�`:�o��eR��������&�ᾪ��Os�*(�m53��(X��g;����c%�!=�md�S:-sZ^񳳲��5&��S�|P�����Ӯ'9.}��^�Hx!���� �~Xnj�m?U0�_�0�%�0�a��&X?f����>7�v��8eſ
j �b�s���ԡS�u�s�N�d3;Y|���z�"�|�'�����A����z��#�xE�6ZaB�Zl',����� 6%O��~.ywc ����5�G��H�5g]�̈́��'np`��=�)�w�n�ʂ�K�F�Ů��>i��Q=��+�rpO��7��I�����˃(�b�e��[�CiPHAT��H�~��s��XY��x\#��xld�lL����!+���B_�P
~��r���H�v��ּW��?.5���b�>�MM�׽�lS�;ԓ{���G��1/�t�}|�aD>�sQ�?2W�:�C���W}���GT���:T�/B���A)���T���V@�Qe�k�����%s+_��
�A8��}������Kv��;�s�n�5}Ѝ>�C���
h�n�� 1�IFߒՎCQĎ���Zs��.��L� ��xfE�R�S�;�M�tX�X���A|���p��b��y�v2��ZK��XF��U�XߡU&U ��i���͔ PS2��'g۰�z�lJIzU_��q��"�Eū�m�ko��H��q5��(PHf�Hr�j�;�Q��{���J	7��J����B��r�������	�MKn.^���;A��pH]"���*���Y[47�,�� 7|���~-���Z�?w���%/�*��t��Q���c�
�vz��/�!����Y��?�ۢW�ub��C����̞�0��/��u֩5��4i�ў?
3&�m���=7 �ư�+����g�ؚ3u�G�>�_�xt�#IW]��z2<mt6S`�^�k�qn>YV����*��ny8|~ˬ�>��fg��o���x��e�61��яQ���'ξ!R�#q	�z$Iw���p�0���J =C�`�����:3�{�C�'}bݫ#����,H-�Ӆz