XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��b妚����Qz9�(x�a��ϟ�f���9p���!o��ߒ(�4D���s�C^ ����]�JН�\�zx���b�q��K;޲�NC]�?�c���m�U� �
;��~��5)� aK���5MGΉRө�y���Ѵz�ϥ��,w�T�;�m)'�?)d8эU.>�Y�9�粍_b�fG�̣ɭܟóN�1�w2�|�} s&u����$m	9aD��B����5����R˸9��ܪ��x��S���.v8��{�,�وL@� Nfq�L��`W�����?�>�^\b4a�/�$чb����:��V5����	F��}�x����X�~���Æ�!٭e�2
a���ahWDd(�m�-��skId�vwaq�e��!` ���?�P�r�b5[�s�L��r~.���ف5C=%Po	�����E����]>��+|yo �,Ơ`�:|�q��<
�{� ���y�^�;���u�ɲ-<�K��(?�a^}��\C�÷���L{w1���/>�����ڝK9{}/jOP@쾪	]�6�=B�i6��
ݤT.�H��BN��rƻ x��՝0^X��'��,5����_5�!�]!MЕ=>�����&�s�!0� s`I��1�K(�`�����g�׹h��Q+f",9�~1�oU��se��1m�-�^�V�1���/r�n��~7�D�ղJh���t��;��sa ���Rdpy<�PvUs�[�����*c���G��g�V�XlxVHYEB    5fea    1830anp4&3	���	 ��t��펑�cZv<
//�H�f�R�� ���%$�eB�f��A7�Si�����B>őh�Q� vk����7y���VS��Á��*	}�;*���>�>&��2�a�Et��|_� �P�W�/��N��v��?Iz$���+�@��/R��lG�N�Ͽ�'��GX�E��6�������F��:�t{n���|G���8������LccE3����D��Vf2
O�:	��e,�M'3��9oFe���,������;�М��V�2��]<@��L����Z�~�r\�.Zg2�]f�H�2�w���a�F~���8
��by�A;Z�`�ٯh3�5��8O�a�z��wM�k}ң�i��������H�)�=���aR�t©�\�ɓ�<��G�f`��ޤ���xm���}H)nI���PA�wx*� ���q�I]�J�:v��c����w���q[^�LͭZ�	cp
��@��&|��
�5ۗ�4������
-�H����m���O�T�p��2�T�����A���-c�xC����\_��rϰ�bݢu�^�
死|D��η0@0鷠�<m��J1AR�=Tj�	�F�J��
��ya�h���i0�s'b ��\4����N�ۇ<�Vbc�-�����u�O�nT	��R�i'T����"���|=�fiT��E��D����4Pa'��Г� y�!�2Y٩jJ��]��᱾S#!�Pc���N����P��3��ː�h��UZ���fH���b\��h�\������2&�=v{��ApJ�>�R{9� �GW�eR(pβ�������}���+p���s!	��I�&K��������H)A��7G�R�A��.�ԥ��u�������ۉ�=#�8��B Ԫ�Ȫؓ�����@�|H���n���Z�t�c�c[W��A��4BZ4��~ @��$/�I @�|B��� �]�P����$�u~Ug�Y������O�X�*�3�ԅG1s��T͋��o���=���șF*>��An��g�.���y}P��o(�:mױL�A�vز����v���BE"1�s����E嘗M�5[G�r"�\ �k����)���I����`���`�J}=>_aI�5�O㓫̛7n�.��u>!�?�Kf8�ﻌ2��C�s��.���:�`~'M��΄�#˦��n��G�Q/� X%���P.M7[:�փ�LԠ��]2�2aa/����P�����(�ȉ���2���y����� \��M{*>��}ݰ��^Lѓӕ�+@[G������zp��wđW3�1��>��/C�����o�o!sJ�� �,m�`�F���k�o�&�N5��nE��p�Q��������u��>�N�Y?��	�Yq�ٟ�<w�L�_q��� V�~�)z� n&���h��� c���5#�4q5�71�=�UXV/ǟݮ^���ؙp��P�ɑ�Q�"n
$T1>�����u��(���$���(
ґ��C3�a�q~Og�4�-���ĹP�����hڧ3��'���Wo����#d���x�lґ�����g�$�'O*&����r�H+�Qͼ�J�˷-��G�|�Q,�d�ɥ��|Ţ~i�R&-HJɖR��N��,�bS����8h�O�l]k�mKoːW�;c(L����R?Kq=��'�I>�1}����j|�ht��~.�ն�R�!�MЖFɐ����K)u�t0α�5��O �n�eιAY�2?#@����@ŤX��-���uf�r�T��"��%s�FD��3�y��fc����} F��,�IYB��g��9�\BGDQ�,�p��`+�����G^a8��3�ق��V��Sk��	�g�"*U�ߤ(��vݞ�6?�>��#S3�1��.N�|^ܷ��` ��������$�:zӱ�	p�"�����0�ZD�ub�m��̓���J�aJ���.�#R�T5g�,�|X�v=�qt0��"8�X_�W����mi˳�[G��Qn�F~�E�5�Ŏ�>��ц�������m;�bET0�۱./]��T3� g�*���4�+TZ=Yj�~?NTR@<B�J@L��.�gD�g����Ԋ��W��^Uqǿb =9.�
��O3�	�{��:kZ<��i"ºx� ��1��[hW=}왒_��@�0�/�!�nG70���ҁ����v�yk5>VMqn6�,��-Y���M�η8d��60�~b�� ���Ok��]P����"z��F5���ޕ�On2������`,:VYBvw����4�5τ��c�/��߿1�-s�P�amj�q�4tq�T���N�h#\�s^�a�]�yev�M��N���n>��@�0�u���|-~=>,���7׬u!n��a�c���Ϝ��v�J�g��t�$q odZ&�sY��}t��В�R�;F���SQ-Ft�}A�0�]�������fn?t%ϕtHp=����C�.�]�9²͙�,xBWQ���3Iջ�o�n�����C5�����k�G�m�`UI�۱ߒ��F5uګA"c��4߱�@��u�^�G�*6`p��8�kg9�Z���o�k���iq���_c�c�`o�6U��+]ѫ׾�����8�ώ+�Ϥ��9x��q�#�<�����)��V�o\�/g��δ�����vGJ�t$��V�j��~h;g~;OW� �	(u��=��ӱ��ajs���do�vě/>(l�i9 ���`�k��<1�����d!��`j１��f�L��BWv�N�����9H!/�/;T����O�y'}�������[���*Ή�Ӻ�Hz��H���o��d��uf�$(Mjo'�&�y�^>��zА�fO�S�"U�H�_�����r�p�)~JQŪ�#����}��Yy���.�ɷ�/Z��5Po"�P��K�=�Xh���s�l'8X}%X���%�;��O>3g�� ݙ��@ ��N�`���U�͉��X>H��%���օ��L�DYe�nBh�A��`m�E)�~#�&D�^�;	Q�O�=�+$�EM���F �OCO$-+{��Y���/�?��ZC��s�o���R�]���Sqsop5I�@;ѽ�Y�㝴ȪJ��}��y=W�"�^��och ���HZ�H��&�l1�D'Y��M�N��ç����K�j�
�l"?`��4���o����f����Hub,���R6�6,D��g���6��b�h�9�"��������s�˃�H`B�]�eH�˲Yn�q�<a��x�J�u�UQg?.0�W�i�fO�u[b
�Q���J'���ݏ���1�z��j)�qH#af*��d��8�p�+Rۺ��.�L��vU����J��w�eW�1Ν�������Y%����"���r[]��� �T/�#5���l�7�������¯��%�MY?k�c��E��R���yW�l���N�ե*��f�v�2�k��Ƶ��u��<)��nV8����央R��x��+�'�7��?^AM�Э��AR�:�6��vR���̫H�s#WPDQ�U���l�p��~�#���[�3�r�e�)�k(ި:@��M�*��,�Gy���e�f���CI�y	�7�KT/�ȗ=�E�_�73wx����Ҋ���`l�W1?����e����$���.˧�Y,x&7ᅨY�2'���R/F�o�Z��'x�+��A=���G>m�p�����1<�`���Lhb�����OFg�?,pF}2fU����. �3\/u{<zN)�(��&�?����j��t��;,%%���r.6W�^�P��?�߁<l:���.UC�#�/!"ǏV�6zf�E=w��D���]��u`�g��T����n_�;E$���65j�ִ�p8��h+^H�1���#�>�O�����C^n�0�MI����a(>�2�9�mۂ	J��f�|�.1�؉���0C�n��0��7ģ�j4�=�O}(1��ޙ�!+�g�0��)�[ƮI�g֍�� Fr��K�{�U��,��W��y���b�y��9����X�ǎ��:�-�9�������F��сӶ�=�f``c�<�'kҢ~4q�]x�	$ =��t=�\,<V^�'�7e��������L�H��>�ᚅ�^�3�V��{�)���4��Z/V�b�>	�+�B�7<p�)����q]+r�~���>ogs���"�Պ��~{�.��/;���`����/��Zd*��s�sz׳�ư&*��b���!TA<�/���=�yA�Z����ANO�5��F�o!�s^!��h����8�͸-�b�R��(��v͐�5�`�.�L2������4H-��n�`N�n�[�K,H�F=U{�	
��a�勔�2��j|�?�0LN=]���J�!�s�$�"�#"}�&,�QϦG\�8e�!��"�C�_������������c�%�k~�I+�[�|W�*�� �W=�M3��mh�+�3��N�*�I���ѩ}� h�[vt�H,ʲj~k��/#�/Sp��}?v���'�e0ײ�x�]�
GT^KT�
���W�9_�8s�}R>���g1�ԡ���K�7��t����̉�\'�dr��l,�"��� ��f��!H�e�,ֺhbf-]M�ϙ����i�t��A�����(���^1G�l*e�f����:�NM�1J��c�b*��O�-��-� ���-x<��0r>O��c�M$�OJ���Ң���h[�z����<Q�b�ì=�dQ��^\�Q; ��	;z8�=k)�,Z�
�V0��y͂�mT�J��u�{oܻ�@Re4���j��T�GL��5�j��2�5ηN'�|���0����a��V'E�� ���~�|�8�֙�P*`$J7�0V��;�>������@��N��kM��;H�>[ʹ����]di�z�o�˻7����T�l��.a�M"	�7b���N{��2����j=pf��\>:�&A�6#.��8���Q$5嗱�-�Dߖp�S�sQ� [�D
�4������Єx�pC�~�$f�ʧ�P��?���r��, ^�b�jܐA��'p�"�����!�����Up��n	]/'�R����QC/�U�*T#DF0�HN�*v��:���3�>	!���d\���+�>��e"��#&�$e�a�f"G"�\VP��ӫ�4����d�<����Xzo�Ѷ3����p�h?�!���3���F{�VU^-��xn�z取���0#��"�|�?NΜ %H���x��h��J�, `�)���񟨷�R\+��a�4h���lRx��ȱe���<��4v��#�u2��L4E�@�v����vi�K�\y�,ȑ�sf�Y-8̀?C�ͪd��)|w��-��ؠO��^v�%����������eh�4��l,�Ds�{���fJ3 �>{u�ԓ8���ݫ}����0~}�r�/�&;��gCP��j� �͝�SlӢ��m�2E���$t3��<{�Vq��u�K�N���ּ%2D28�ZŇK�A4_cE�g��j�ã�z�@���� ��[(����e�A��
�TV��R6k �s`ŰwF�Ӓ~\����n!���ﴂ����3�ToW��솗�Uǥq�xWB�R�-)���%іm���!}�����������؏p�h}?~�o����X}�G���� �n�[�k�J����w��BRT�N��.*��,WG���[�:���Oj�6�3;�,��y}� �q���lλ�8c t\NxC�4��q�����=r��6k�{���ǒ�|�?D%��1nwJ��O�#�E�Ø+��w ���j3��~�ƴ����[T���
�بZ����4D�-n��N�N<���Y�!ܕ�K�U"T��|x�h�5	2�ͧ�$�8ڜY�r2�':��-v��Vk�Q���[p/����~�&&�ѩӖ��b
�_�� 7(<�Jj?9�T��q��������y�]��Ӱ\���5�yQ���eԨb z4 V��Vƺ��bu��X��m�\�S�@]���