XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����������q TjIY�]��3�Z�iX[k�4CB���k�b%Bi���W\�HAS!=��c�J	%����U�}o<J6r/<�!�!$���:n��i�f�$���bn7�~�v/5�O��uq"^���[l�pdٌ��fl�b����+Pa��P'�@��P����`�7+<99g9�=��%�mi"�N�x���MݖQ�,�J�8F�ui�;m�G���k�.~]`���P������=�/��\G���z�tG���u����p�'J�)>��W�p3���o"���Of��D\[��&�jm��i�)ED�-o߮���W a�cn٨�%e��(�t�[��f��O
_C�,�1�������zC���~
�lE.4��W'U�ڍ �g/�_��86���� ��(.����@8�W�~�֬Q�\f2|O�/��L?V�����G� Ip�{Ȅ�b�3���-N���?5�ډ��d���6Qݸ�;���v��$�9s�Qԅ@��Ȭ>�,�7������A�@�(B��֡������c[+�Β&H�C��+$�	�N���;f�QB��x�wfa��v��f7-��ɑ�ڽqH�,��V��7�\�ʻ�cq��(B'�)�I�Uϑ3�Y��<{Ϧ��}�`#o���,���C�f�P&U%�6���fh�6��$Z�)us��n����L�'ć\��C��|X��Y�p�3�i��/ �!ui�&�h� #�V��q!�M������"�^�k-�Ci�aMF*XlxVHYEB    5e2b    1530��%[��euz�aI��- %��/�������N.\�VEp;
�d\J�d���&8)e�q<��ͳ���=�����:d���Κ� ���˝ώ��)] "�/b�d$��)ߵ�K����ؒ�*�W��Q�ygJ�q�����Ig޶�^ń�wX����Jj]r��[3����'� O*w-y��:pCr�%Lp?d�O0�]L��O��֓��bmܞh�F�%V�U��=oY=`7�כoĊ���YL���@U��I��PH�����w$�Q���+����3���ͻ�7n��\��ri����j[5ſ��?���v>o�h���N���3�m8Zl�ߌIF�|N�o�� g$��7�Q������ld�F{q�n��#�pbX�W Ҭ�Rg����p����`.ꯏg(f���u2|����_���Sӎ� ����t�q��Q�CT�W�nP�˲tI������&m\�wyL�u�+")�Ѭ�,hN��E;�(��*ត���M*���g�ێ�~�1B��$��oI�]l�ۥg�.���A�zٗ_ ������ ��?�^u�'&�{�>m�_Y�z��c�EhS�C����4:��������-�5�R<ɼ�-�P��*
)��ޏC��^f�Ú0��1X��b[���/*�%�X�K�8��<�]�s��lP�uB�n�f�?��O#������ݒ��e�18�ꅤ9(6H����7�i�oփA�Iʃ;ZVËT��2R��x�.`A��N�\ٶ������܅�]��u&��c�k����*�vԚ�$"h�l�t2 @���s��1�s{lkV�h'`�8��'��v.���F%l�Ɍ������?Izsc9��y�x��6 "'���!�!Ӂ^K�$�,���	��Ph�rӻ�3�٠ݒ7��&<�|I���:�qt����g�����OK{�3�V	������=�������i(Ap���z���k�%@��뭖���$h
v掔����p5�#��!I��{�.$��.�v�XG�w�IsHwz�:�)�Z�sGS&��jok\�Av������*�mWr9�Őhr�Qn6B2�M~�S�|a'�_{%�X8��;�;u�q�k��;��ZÒx8%y�zO�7;�*�����:˰:��:�R����GQ�j ��f�xD��:�[�ȞY�4�'	��2|<}P^W�=wdEyv��ľ��u�%�_T�:X�-V����a��
 �\��&?޾�ѯ�
q��(�﯅�zl%�|�(�a�Q*�\�U~��8���o��e'�`���L,$Y �/ƅ$Κ��
�P��6�W��:S���RT�7���^
.���������{/UF���RLGy�bQ�����y��ӎ8(�4��5���%ҿ����] �����A�dY��e�gbK���>ː���T��"@=>:�v�E�"��M���C��-�&i�r s�	�	��ŭ�y�n%��wc$�4o��֤&J�h?��#]����'�B*BK�GYU��S7�c����xJ��?9�[X�w-ߦF�0��H�E[׎����p�'p`��t2D�����<�o�*3�I�h��Ǉʖ3q�\;��#_b�8��j�<2���N��>�^,����HA|�͒e��W3�w�����d�^�_%����r����/G���@��&�D�Fd݂�)���Y��8sGrJ����p	E@��dC��l3�@�1֓(P?���k���hA�QIH�v�ؒt�KYg�Ǜu����ϭ�Z9A�������F� iΥ��5j���y�R�13�C�N�89��M5J�<i��.儙.�t����E�#��vT"��52��^�� �j@�C����*���U�q@B?�9�}f�?�>�rbe���0O>���c�1!������2�{�I�D�R���V�w.݌B��y�FS0�Ǉ���rЂ��T/y�O����-���v-Ϫ�������i�K��T��^�#`�悻&	�M�1��x^d\9�v�"*��8~��k�+��Qn���M�h�C�����T��mY����sU���V`!]Z�Q�FO��֥ܭ.4��ޡ1VCp�\M���/�vW]�5�vh���4M�cK|�y��?;=h�}���]�z�O��"�1G�J�m�5���B��SW��Dc6 H�]q�k�\�y[��H�Αl`>�/�A*��~��Ņ9�9�ɥ�j��َ����Z=�(�R�!xn"jP,2l�7�~9&Tҵ~�������ܒ:~�z�5�+q��y9g�F?�����[G��h�`ə�I���d�t��Q*r����g(�����������Qװx���Y�;�<��w���Ƙ� (W�g�	�~	�Z��u��f��dC��e�p۝e��G=
�O�sD�Xܑ�h��_��
��kG4{�����m��4�V���qE�:ණ/??{��H�3AG=@�wD�g��#70���Z~�u[�g�DPZ���h�jMn�wC�4ź��s��1����+��T�r���Ti�`��_qbU,���jq���cɢ�4�)���ċ���m��Z!0���^\��0��7@7ҩ�I��/����dKY���K�4�O(�q�[��g�b� �����Iґ+��'�TM]�&��'�J�Z%z.����!T$�*�k���]O�N�s���65�k_��������#=O�ik�?�K<���F�4�̂��b��O��˛\D�+��5���g�ů0ET�X�T�2�Ĝ���P$l�b�bk�p'�����I�]g<H����J�e�#�(�0e�}���c�!��Q�7TAM��)�ux ��M	\�)p���=l_�v��L�jL%V�ͺ_���劉�b�&}d�&����ґ㜣�o�3QX��g�n���v�|Q0t�=]ղ�4�1QG��BW��ߴ	��'������ڥ���x����"�}}g�-��!��G.��U�.��l���z����{����揎������ n�i�-����(y����g�I%_D@�˓�� ���&wM�@�	A�nqt (�(�پu�C�>1��2�c�"�c�{�==ޤ�W�j��7���etx��$_��<�A�Qg�����>rWB��f�r��2?�:� ��]�<�#N��#VQ7�����'��@J(n�p����f�5oN���l\���]Y�]R�.�s)�� �ՙ�v��
LIK'�YK�_tī)��o{L�@eE_�
�� ���RLo��É2��m��j1��S�7���Tx��$/+,�fM��S"�Ƴ��>3�)°^p*/�K!J�LH����� ���P��t�3H����z�:���97�f�u0��xM��֦�3?���w���M�O��5�W�	�&��{��ڜ�
F_�
J16�Yk�iniJ��1cQ�>��Pa&�`<��]���yO��ϧ|�EP z� S���9o�x���
	�Sڇ��x!�LL���WNcuM5��Tx���EG?S��\��
�C#EGT{�?l�Z���$�%���L��}k�se���b�pQ֫	�ee�V�V֍����;g���Kn";꯷��^��>ۛ��\�?����� ���S~���o�B�1ϭ�1���s-���bf�jg�RO�����}g	�ee@V�=f�������[����n��hP�_�ˤ�^>���|�}��)�vy�k̈́�|�32�y��&.Ao�ֽc�����^�6�Ｎ���*}����Q?���L�m=�E�0���������n;�Q�`L�]��6�L�.ȴ�\d�Y������X8`u_<�i��|�=���'���Z�9��u�ҙJ9���+�`����1� h�,-�@!���Uv��g>Oȗf3��-dy*�Ɠ������{��޼v'�.o��;*"e*�cS:�@O���V�-ۡ��T��[k��|<"$g�;Yb����(��Kv��T���(e
���f��ddJ��2H�����<4i�s��O:�9�?�ѦP��������)G���!P�u��ǰl�:��F!�G���@{?U>
,�����r7ߞ�_�="\z������"QS�14�葼��]O��8	���&.�3C4&x�xxi��;H"E�L������¨C��6�ǟRӓ�(���z�P�Q�!
��lpΤ��D+J���8�ju{d��>��ԏ��UDDj0�,���&�3��?F��[
W���rG�?�%�y��#~�6��M2��\�w��)�C	�P낫�;���Xe�T�DF�o�ٿ���_+��5X���|�+���J���#i��"9��7���"���R�M��v�s��Gy����e"���AƖ �VmЇ֡48�Q
�ѐ�#ï���!���aޱl�9�A\L*!�H���_'�e	F��]�q�!��hv�o�t���Z�6_��HG���?�]<��zU8��Lk�E�s�T �,GERύ�'F7\��6a��ViW��L�H�na
�7�W�-I#�
�e�vN>��>�".�ɋ��K�(��%��++�6��T��ߺ�GU�� ����w����~���p�
!Dh~�g�}nY�!n�}pv@�@��r��S'P��}�|��ᓀ.+�9X�vh� V5o�8����m.��h
�	o�s�(U��&(B��*�AH� ��MF��K �93W���s����S�#z"2�̹Pt�+��#�R�F��%ωM훅F�#�=�W�-p��2NP/�6�4P��ヺO<o	r-���uj�$y�X�[Yߙ�Й��u���8d	q��	�����P�ķ�,]F���F�^��!/�$z�ͳ�g�צ�2Aצ%��f�����7ce��X�ƍ��pd�����!
�Sj�!�B?�b�l���_�	�n�!Q9{ekλ�mȯ�]�U� q�j5t��ښ��s���RϪ��r������4"��/�r_���M!�>�$�R���C�J1��hE)�T��)�}��3(� �%~l͎G��$�ͨ��acN��@#�v�=%�^�a��i��L\�z2]�jF�}�,��[?���s~�C���9s�R5���dX����|�D��D��'���Uj��h��ƒ���1ꞫKW2�f���Oݜ��Rl^�{�6_�=(��N�y�2�_�2T]�n�)i�PE�ڙ�"O,���x�2�{p��~��H"g���Q����q��\��JN���z���۞����kګ¶���%K�9J�xp1�Xc�����3ڜ���2GKd��}6�y��}���T.O>