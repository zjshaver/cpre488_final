XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���R%.��shA�K�������R����u ��b��,�)S���p�@�(Ӕ��%D��CaW�}f�6	�2����.���Õ&|� z���� ���B]�<�Rl(���^���Lѹ�J��*�"��T}0�4N �f�U�� ;/`�t���8C�G�Z%�w�G1����j�~p�vp����"�Z�ZMK����$c/���,33ԣ2�=�3���9�������H��$�W��	dl�]��I�?��-��ǋγ������j6��V����.��y�J�!�� �Z>s�@im��>_PKr��I��z���h��|8�J���;��4����7�S���:��3Xy�ɩNKJ;�J���&�M���h�F;E���Sv�p��=K�5̝H���E8�}yʖԋ-��ߜ
di�Q�=RLV����O�Ms����w�ّ��A�gu��_~�Q��(]��g���A�U��ɫ��c�+�a,z��9�a��Q�`h%N��õh�t-WX]����*xO�ѝh�=�:[Tx�v[[n����W@g�G�O�nA��
p��� � ����N�b-?�Kb��[�%�C�<��e9璠U+i��ǉ��0mۃ�we����0��d������ti���0�u���l��1���i.P�UM����A~���4�/�4�?*�r�P-�<���]�,��_߄䛨+��Z0+���������U+�<���jV=�V6����}�]=�����	%�UXlxVHYEB    5d29    1390ׁJ�H�B'��ߢq� ���Ѻ���j|S��m��J�4������@f�?��^7�6�O�+X��9n��O� ��<�G�!p�Zv(|��n�(�mՆ�Ɗ����W�'�_J��<�;�z M�̖�����w���ȵ,�v������!�\^tz�(t^�7OY#V	1���#O�0"��{�'�R`l�_
��h<lD�>3�e��y���ʩ��d!�9��q��Is����XB��5���RIo��T�ks����Ư�Jb~��q���yqmUm-�R�	�˯)M��jS�7&h�Q١�j5@M뿊�{Q@,�D�3�b����Ѳ�D�=`��?y�R9��ROZ�N�RFQn�g�jY_[%�r��s�jc���{�F��.��&"�%�G��
����`KřIbz{*���ˢLC��b���̨YEy�CW�~���n��Q2�I��H9���Ŭ^G����1����Pڔ��d2GX2T��ԉ3�T���<zmm8G�%�f�g-�;��F������Rt�p������7b���Ʌ�B�@�H2�s��NL����sml-O�� ��~�=�9į����P%d$u/@���%�
%�Ed�K��n�.��V�eK�#�c3H_w�O�^�w�D��nb��A����T�(�j�S��B0�Dd ��h��ۂQ:V�M
�d�΀q��r	*{k�ϓ��%��� �.���ƁjE����u�	x@իͼ�5�񵬬/��`mt^��pE���d#؀4���[�)�dǨ�
���\l�m�#��w��y���qf�7��\(BE�w��:/��em,�=C���k{����c^�M�+uS$�QD����&��;������� i�oD�ۡu�ߧ�C���=��-��\V�T� P�t�b�xU�w0���E)�5�<G��B1Dg�l)u��]����n���jiJ�Q&�o(NY`z�&�F
�ߐĕ�a�[�hP�b��L	0�41��c<Q����W���Q&��%���;�E�՛���J��)�cN}��4��������b��tys���8%^��en���8�C��b�@�o�z2�+�ߡ�v�^�#* i�9{�B�ɩ���UzU块r�b�ߗ"�6]�����!�4�����YQ��E�$�� }��	���!	 M��t<~��j�_<_��2��҂��SCN����r~� =
$�}�qH�.q����>Mޑ0Lj��r��<�E=��Ϗ�`�q��KT��1�Q`����=��2��.v�E)h#��#(�>D�caV\��#L^g���&^`���t�
���2Y��ZW��X�xC։-~��@ �.~R��9��{�1���k�4F/ۦP󿉿޳?�Ը�f�̺�f4ܜ�fC{a�1�0���Ɵ�� m]e���ֲ�ëb�s,��!"�8�����|#��*=�=Yv���>��jdF�5w�����V�⾛e|��iFKH�H!ywV���5j#�sS>��rI�wʵy��@FM����@lT�s�'p���t�f� ��U�@F)&߾7,��yR �J��Ж��I+���E�h��a_��K�(A5��q��9t���A�!V�(ֿ�1z��o�C��`�z��P�y���4j- ��g<Ջ9����Cy�*b�
�~��d�6���Y%sx}
s�-}�q��4nM~�J`��j������7�{K*�X^�{!b~���ޭ�� �+.0]�<�΢u-/�<���z�x{̉��T4g@���ę �4U��(w��Ua��+�V�@�-�Mֿ໎���Ht?�
�U�T��N����1Kb��Ip�h~<���Ec?L�WxIMW�������gk��H��_���$Xs?N���ă!2#<���#D�h[/q͞�S'��6s�ۮ��Hm�2
QϳB..xߪ�"�F ���S�r�-=�U	]������yM�����ނ�q?.˘7��yࣅ��dsv�Y"���mB�e�'��%6����샐��Z�Hy��Q���PJ�h��M�~F�(�����������.Z��ZG�!P���s��g���1¯n��D�_S����"&W{�v�A�ioY_�I�����h���F�voDAB9q�y�2��wP���v[�:�;c�s(L
�(�.�lѾШ�w0��f��#78�a&*V�N=��G�aw����m�
gI��'9��k���cW��,%��muN��v��S}LxuY��\#{�Q�K�X}*�D=h�pL-����]r4 �*����v��3rR6�\�OS)u��)S���F��cMH�Q8����T��P!��n�rըW��УoB@*ǽl[�	���
0C�l5��,qF?r`����p��ċ�݆�Oɛ���D���N6yMвś�ܑ�:!t�S�u��r\�l�g/13�ހj�6���B�|��f��a�};�n�6d�[�e_����X�_��3.��R�����	�XgUp�m׊W�!��F1�i����v�*zH������1>h�L�!&��n%Ĥ� ��0I��T��Ez�Ġ�˃�@�B�pr"d�[�.0��i���I��e�R�|a�}���Ҕ���7�AmߝԢL�v8U��gW����j�I�!���)�ى��A@/Ӛ<R_DW��PC�{�d�N:?)(����&�hy�G��*��^kC�7L����,���s` ����g I|�s�(c�p5���o��C�[,�ţ�nz;�����.���Ǟ2)���:PC��O�x_����vLV�go$��1x�x��>R#�J*@���Tس�6~���<%�����r�b�y)�v��\���������ֈ��ڌA��`P�5ag��N�M����K��`�o��0_���n/K1Ln�:= �=�jY��к�)�6���(Ԅ��KY���6��x	��a'˷8�g��������z;�  �\-�V�ϣ#�,�ށ7G]���l��_���L�;�&�x_a=T@[S��fE
K������e^KH����I\�(�����gڍ@)&��mfI�j�v�ۚ�?S"�Y6���\%���h�h���{0�ym��L�)��T6`�������b`�~X��惦������lq}���/|���~vW�@��N|V�ؿ�͍ӿQ�c6�Z}�����q6����"x{��({����-?�}v`��ڐ:�W��MJ|�A�Z+���q5��*<�bH�x�����?�a�bA�¨�)�|��t�1����xt�E�騬n��ex�#�
]��Ƌ�}�z.	��^Q�.Ya��m��Bk�s�*o):"�蔼��d;ͺܛXs�>7�'z�_ZI>v���^kF}�=�5�h
쯯�IS����4�:4�4P6��ұ�j��o�9����<g%`���W��YM���O��8������!��F41¥5��`@��>5�V�@/������wB�T��C����!j7�\0��ڔ���5��9��7�� ����a舜�)/�����3��g��}��'�u@uϸ�tAjՋ��R�fګ���_8�g[����c�Ӻ-?5���Yw��Ao����F� S`%�2�"�ŭ$&<���������� !wAf߮?��Y�`�;#U�J0.q�������C/���B��@#;�3����M4��u���3s��@�i���`V.j=�?.��f�#I�T�W�t��,�v1�{ؒ�g?{H�F�[�
��M�uz@�t�E�=]m��Oh��{2Q*!G�	��eu��I>�j��i�ph����QЋ���f�+J01j�0���p]\GXS��_Kt�3��}���E,A�+,�5�����ZO^�l�$HU������b������#����z��n�ż�F�0�a��ö��%qTwQ��#f}fÞ�b)���/V��F�=��5��S%�L�[�5�����/2��ގ+�bA��a_�1�<��G�^�D���%5J�1+��-�#.�_��=+����������/�b�ѧ�����l${�3n�az�|�v?8�s(\���u�.{�8	m�z�����K�7a#��\�ney���e�$sa���}�U����F;���y�B@�o`�0@�!��Ѻ� ��B�B������)�v���G� �"YE=O��'�j��3B��ìZ�!�^�!���x)��0E�~���W���W�p�rl-�JeuYy	x�(VڇD�l��m:/j�`�OQѧ:}���3k��V�<���M�
z���T5?�↝>�r4t�r��1����� t٩���K!��?U���آ]Y����u�F����?r0��N$#���L�Z��,���#q+O;
�1A��S��cڸM�lVѥx!Ld��3�p�!8_�Lp+�i��C8w1N1L�突if� ���bC|b9�8��fV��1��]�'ɹ6Zx�~��s��&Ruw<'�U�zNi%ܷ���v(J��T�S�:v��B�����/O2ψ� ��^[��`I`��Mc�ր.�q\Fd�r?�o��7,͎ �T�Q���|�9�k���ß-^��9��+����.8�)�)��u�_�Y���>��Y��G�q�]�5����}C- �pSmdό�ޘlP���H!�:�j���qs��V�K^�˻T8"� ���*��5ڱM�)�.�4/%j}Bd�J�R` ������*uG)�b �<iɀ��B̏n�WP��7v~��U�P9Oٰ���Uҹ�{�<�{���rU"��H9g��P|��r��0ݼ�5#*(#��<yF �X���zY��l��@+�'�}�������V�[�"�U?�N@�bl��y��vmN:�$�c`��azw=w3$�[с���[1������*�2��7���E[��