XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��)��cCl� ��<�脴�QR��BS�(QJZ�u�t3H!�{(Ax�>���3P#d ��r�*�ZE�h�B_���P��}��Tt��#���f7k
��+��S�KT����R'�`ˬ�JTY��Q��*�U�*��gq�?-�\��<�o�9~p�z32��)d����j߹0�5Wd�7�t��8W/��9�ߨx���n��Z�VBH��I���V�b�(�#�������5UU:��e�}�h:<�ҁ�CT�N
��E��0l�6�_���v�n���"�aO�NI�d�����"���*>�R���ZW�Ƀ���YaTU.�gMJ�HuLҰ�ԏDh�;.gWU��A_��|��x4�з�Z�� �1#ڤ\s�7�7�p���(��C��n���]M/G��P����Z�����
�+m�;%�d*� �lD��y3��D�}u�`�>H`^���L�U��Օ��)�gì��0<ˢh@n�aƺ�J���@K���1��7V0��+�,��ؗ�����0xG���d�Jf�^�8��xAbK*��	پG�p�.�N�js�ࡹH�(��д0<rH�.T�W�8�Eޔ���K;�/�f�����^�}z5������f����xG6��Oc>�|N�ħmS��O��׻^��Hk�u��|��Hy�#u��Пw�f�
V�0~��
R9��8\v�c�{�-��`
�������A��xy���])�)zJ��տ?� %I�e��z�H+��6�<XlxVHYEB    3d1e     fa0��BQ
AMaNJ8t+��b�g��z���'>�/5Nf��;�-̓�D'[�N@��D����n�8�~,jO�t���d�]������[�%0P%�=t�"y&|�v����P�d���	�����YV�����xG)7B����i�����[;7�9�Z�K�Ӏ�c:����A_�
�|��d�2#_�r�1���_x��f��,�7yFŲ^�	Ag��/Y$��Q���3ڻ��h���0.*�ɺm�}���!>?�͇�uDO'��T$�a1bd��6�)�����"ͭ��w��m0m��kN�n�q5 W�n�ɟ�zu0t?W� M'������/ ��6�$��2��^�ٙ�u��佢R�	�^�1���+�8�:�#dK��&����N�b�n�Ĭ����Gи�
F.�>�7K����4%<�u4;N��@��ؖh�x����o`%�'8�گ�\��%����
��?�v�!x�6d���!�\G���M{y1�OM"���r�YV�8K��!~�Z��U7"�5��sydKGHKؠ�C�O�	.��?*#D�Gx*-k��`��<�(�.W��T��&r���&|��HT��g|�)s⚛���9Ln��	l�F�oժ���[�<�O�Q�����Xk�J�a)׽�����L�fO �^2Ł���
"A	����V�͐,�K�J�/�j-ɘ0 ���ytQ�`��޾T�����t#��f��#L�{�gĲ24��p�[�Y����و�\�aDѫq��X^��~��rr�h&�r�8�4y써 ��la�����%�,@�D�z�c 3�S�K╴#�5���g�{-�{��Q��%-5���q77�QҼ��ml/6u�?�XQ6G<b0-Ւ�t�)a̢�ϝc=�"��@.G��UR2�S#o ��w���X��i�|���C�Ba��"�L���x��ն&��A�ר�o ��^8��`?F���X�e�(����+&8
����ǀ �_"g�tl�OE~N��Ń���N�W��5�k[��e�(2�fqѾ���si��Rt�W����A������<:�uk> N�j�mg!o*T�YOa!�� �~A�ɱ�X�,3,1���:B�ܰ�,�'��@��8(��>�}�������<
�
��621FƎ������Z"U6�a0�?� �;���߿���B�͊	�ݶ~�ت��,
�3�*v�$W���䪄��D�q;��2��r{B���.DѠy�8v҈����Zǒ(���r��F=>�n.��)�:NM�	'p�Tf�٢&���� gD���?}��Wc&`���s4����z��5|V�>�\�teb1���(��	���6�/�.��gdb/�������
Ͼ"r
���>�MT<�7�J�GB�0�1�ͭ4	
���7��x!�J�1${Q�G��"�R:�Y9�]���)������e#���3� \~� f�ՋX��E"������u�6=;E^qԒjI5��x��pfTD�ˠZC��f/�s,f*j��"ox�����g��oLQb��F���'�n⨦��j�t��ˣ����_�A�4 H��7��(���G^��K�z�Uj���|�u���z��`�g���Km��%�Z�*�#*�����*ǹzr|p�$���B{|D��^v�j�B_����f��=;�w�whP0�U�\,��"�=���o2��!҃�#�o{a�_tCU&����3a{����tPW�F$ź��,%��J���V���gOp�:.�*6Ƃ۬�P�XY��r���b��ۭK��rZ���&����6��W,���K�<-��ͮ%;Y��ǌ�!d0ġ���ȡ/�e�u��@��r7�����s�8�6EC�\�6! �p��+`'�f��@���h����GuX��e!:�Mk���a6ҙI$=�+��4_�B�ܼ����a�<n�P�5�n�Rw��#�/I;����&�|�� q��,��7��ⵇ:��ԆG���y�!!�!���
A��r3���l�"5�|h���߀���n,�O��dȫ����g����~��ţ���4��rN�(�P�����O�q�zd��*ԡ$�!��3�]�����/�Wޏ���Z�G��#��V�Dà���\�h�K��$C���f��A��N�@�5��/�K�l����Y{����7n�E�e��ğ���p�5 wv��ck
f]��0�~������6��-�n�9���ঘ��¥jh�G��6�o�ā���v(��7��j���c�^x	�V�pOT�Fks�m��˂����zgc4E��6oSF!2 (:3#9Mֱ�4�)���9���#L�w_�(�N�&&i��26����f�Q����M����'��E!ު�G��W�Q�{�cx6�.8�~��)���dF|����Mt��a�ڲ[@����jS��y7�pj:&(ğ7>?yR{��)�_���*�gha߅�W9�G%N�az3����p������t0���/���rik�EM�a�n�S+���@�CIz�*��	'��K�#~�c� >�f�a~i��D�D�Wz� 8�=�5:M�Tr�A�$0�1׆�n��5��²�e�����r���l�:[w*������򹇻��jS�6�ӂ��T{稨e�B	�e�р��TV�}P�����]	��0�l1�=�����_�|�do���@Wd�KZە�8�?=�{�,=�~��CK��ܩ�-
� �:�I���@�����-0;D.�j��5Aa��F�����0�	x˩!�-m��s�d��yF���z�����m�zk��rj���1L&v�ӷ�"���C�b��������ݥ}���/[.U��;��o-���2�����XlGz'M�8�:|���7O���ӥ#�x7�%�2q��n��?��3�n��uT؄!��)��X���<���	H�d�E��M�n�5�9����n�K�A����k=�6�sպ�$�.9LO�?n1eQ~��v����k*�Lz$p������;�gN�����k70���DS8�@�]�����#�3r�P=��K֚;����^�n�tJ����z�^fP9Ҥ}́��y�:P9v��r�zv�~��I,�-���3]/0�h=�B��׀hނB�*�bˈ<���<��>�i�p�q�sV)f�5��X���٭��ޗ�"�yC������/1׻a8o<9��gCN��|�|��;�i��d�ET�fM!\���휷�Of�c:�	ߊd��pq���_��=T� ʢ{=C�( ��I	���5V�#lzǘ�Nd�v��^����s`� ����c�9�2�W����#�A�%Q�|�����1�AkN�y��f����[�΄��:\���n�A�~�Ae���ns�c"Y���!xj �sN�~.&���w�3M<c=-��.1�M��຿�>��F*�3« V+Y�������D�Ϡ�U�EU��Rɭk�O��u�4�`<���aHOM�����<�"bw�l���U4�r�2ՂG��\7ұ�^oS� �p����5��TdN�NH_� 2�-}?n;��0�nn�&5n�|P(����jT��?)�"hX��g����ޭ6��i/L�V�ZZf�y�`2V_aJ��>���I>���bĩ��^W�a�'��(n+m��	���l�w,�;�8R��s�=��=q���t������|8�L��k�Slo��B(�f�`S<BB[<ҧ�a{�@�0"u�]0f�A��A�3��6��SƝ���u��z!?W��KVC�A0�c�c�'����-mUD!����k��s��8������	�D��B���YV�h�$�O} 8��v	O�����F���_Ep}�9�9��׿l��G�%k�s)�do��Vyv>H���)��������